module rotation_factor_4096(
    input                             clk,
    input           [9:0]             k,
    input           [2:0]             stage,
    output    reg signed[15:0]        x1_re,
    output    reg signed[15:0]        x1_im,
    output    reg signed[15:0]        x2_re,
    output    reg signed[15:0]        x2_im,
    output    reg signed[15:0]        x3_re,
    output    reg signed[15:0]        x3_im,
    output    reg signed[15:0]        x4_re,
    output    reg signed[15:0]        x4_im,
    output    reg signed[15:0]        x5_re,
    output    reg signed[15:0]        x5_im,
    output    reg signed[15:0]        x6_re,
    output    reg signed[15:0]        x6_im,
    output    reg signed[15:0]        x7_re,
    output    reg signed[15:0]        x7_im
);
    //旋转因子以2^14量化
    wire            [11:0]        address1;
    wire            [11:0]        address2;
    wire            [11:0]        address3;
    wire            [11:0]        address4;
    wire            [11:0]        address5;
    wire            [11:0]        address6;
    wire            [11:0]        address7;


    wire             [9:0]        weight         [3:0];
    
    assign weight[0] =10'b100_000_000_0; 
    assign weight[1] =10'b000_100_000_0; 
    assign weight[2] =10'b000_000_100_0;
    assign weight[3] =10'b000_000_000_1; 

    assign address1 = k*weight[stage];
    assign address2 = k*weight[stage]*2;
    assign address3 = k*weight[stage]*3;
    assign address4 = k*weight[stage]*4;
    assign address5 = k*weight[stage]*5;
    assign address6 = k*weight[stage]*6;
    assign address7 = k*weight[stage]*7;

    wire [31:0]x[4095:0];
assign x[   0]= 32'b01000000000000000000000000000000;
assign x[   1]= 32'b00111111111111111111111111100111;
assign x[   2]= 32'b00111111111111111111111111001110;
assign x[   3]= 32'b00111111111111111111111110110101;
assign x[   4]= 32'b00111111111111111111111110011011;
assign x[   5]= 32'b00111111111111111111111110000010;
assign x[   6]= 32'b00111111111111111111111101101001;
assign x[   7]= 32'b00111111111111111111111101010000;
assign x[   8]= 32'b00111111111111101111111100110111;
assign x[   9]= 32'b00111111111111101111111100011110;
assign x[  10]= 32'b00111111111111101111111100000101;
assign x[  11]= 32'b00111111111111011111111011101100;
assign x[  12]= 32'b00111111111111011111111011010010;
assign x[  13]= 32'b00111111111111001111111010111001;
assign x[  14]= 32'b00111111111111001111111010100000;
assign x[  15]= 32'b00111111111110111111111010000111;
assign x[  16]= 32'b00111111111110111111111001101110;
assign x[  17]= 32'b00111111111110101111111001010101;
assign x[  18]= 32'b00111111111110011111111000111100;
assign x[  19]= 32'b00111111111110011111111000100011;
assign x[  20]= 32'b00111111111110001111111000001001;
assign x[  21]= 32'b00111111111101111111110111110000;
assign x[  22]= 32'b00111111111101101111110111010111;
assign x[  23]= 32'b00111111111101011111110110111110;
assign x[  24]= 32'b00111111111101001111110110100101;
assign x[  25]= 32'b00111111111100111111110110001100;
assign x[  26]= 32'b00111111111100101111110101110011;
assign x[  27]= 32'b00111111111100011111110101011010;
assign x[  28]= 32'b00111111111100001111110101000000;
assign x[  29]= 32'b00111111111011111111110100100111;
assign x[  30]= 32'b00111111111011101111110100001110;
assign x[  31]= 32'b00111111111011011111110011110101;
assign x[  32]= 32'b00111111111011001111110011011100;
assign x[  33]= 32'b00111111111010111111110011000011;
assign x[  34]= 32'b00111111111010011111110010101010;
assign x[  35]= 32'b00111111111010001111110010010001;
assign x[  36]= 32'b00111111111001111111110001111000;
assign x[  37]= 32'b00111111111001011111110001011111;
assign x[  38]= 32'b00111111111001001111110001000101;
assign x[  39]= 32'b00111111111000101111110000101100;
assign x[  40]= 32'b00111111111000011111110000010011;
assign x[  41]= 32'b00111111110111111111101111111010;
assign x[  42]= 32'b00111111110111101111101111100001;
assign x[  43]= 32'b00111111110111001111101111001000;
assign x[  44]= 32'b00111111110110101111101110101111;
assign x[  45]= 32'b00111111110110001111101110010110;
assign x[  46]= 32'b00111111110101111111101101111101;
assign x[  47]= 32'b00111111110101011111101101100100;
assign x[  48]= 32'b00111111110100111111101101001011;
assign x[  49]= 32'b00111111110100011111101100110010;
assign x[  50]= 32'b00111111110011111111101100011001;
assign x[  51]= 32'b00111111110011011111101100000000;
assign x[  52]= 32'b00111111110010111111101011100110;
assign x[  53]= 32'b00111111110010011111101011001101;
assign x[  54]= 32'b00111111110001111111101010110100;
assign x[  55]= 32'b00111111110001011111101010011011;
assign x[  56]= 32'b00111111110000111111101010000010;
assign x[  57]= 32'b00111111110000011111101001101001;
assign x[  58]= 32'b00111111101111111111101001010000;
assign x[  59]= 32'b00111111101111001111101000110111;
assign x[  60]= 32'b00111111101110101111101000011110;
assign x[  61]= 32'b00111111101110001111101000000101;
assign x[  62]= 32'b00111111101101011111100111101100;
assign x[  63]= 32'b00111111101100111111100111010011;
assign x[  64]= 32'b00111111101100011111100110111010;
assign x[  65]= 32'b00111111101011101111100110100001;
assign x[  66]= 32'b00111111101011001111100110001000;
assign x[  67]= 32'b00111111101010011111100101101111;
assign x[  68]= 32'b00111111101001101111100101010110;
assign x[  69]= 32'b00111111101001001111100100111101;
assign x[  70]= 32'b00111111101000011111100100100100;
assign x[  71]= 32'b00111111100111101111100100001011;
assign x[  72]= 32'b00111111100111001111100011110010;
assign x[  73]= 32'b00111111100110011111100011011001;
assign x[  74]= 32'b00111111100101101111100011000000;
assign x[  75]= 32'b00111111100100111111100010100111;
assign x[  76]= 32'b00111111100100001111100010001110;
assign x[  77]= 32'b00111111100011011111100001110101;
assign x[  78]= 32'b00111111100010101111100001011100;
assign x[  79]= 32'b00111111100001111111100001000011;
assign x[  80]= 32'b00111111100001001111100000101010;
assign x[  81]= 32'b00111111100000011111100000010001;
assign x[  82]= 32'b00111111011111101111011111111001;
assign x[  83]= 32'b00111111011110111111011111100000;
assign x[  84]= 32'b00111111011110001111011111000111;
assign x[  85]= 32'b00111111011101001111011110101110;
assign x[  86]= 32'b00111111011100011111011110010101;
assign x[  87]= 32'b00111111011011101111011101111100;
assign x[  88]= 32'b00111111011010101111011101100011;
assign x[  89]= 32'b00111111011001111111011101001010;
assign x[  90]= 32'b00111111011001001111011100110001;
assign x[  91]= 32'b00111111011000001111011100011000;
assign x[  92]= 32'b00111111010111011111011011111111;
assign x[  93]= 32'b00111111010110011111011011100111;
assign x[  94]= 32'b00111111010101011111011011001110;
assign x[  95]= 32'b00111111010100101111011010110101;
assign x[  96]= 32'b00111111010011101111011010011100;
assign x[  97]= 32'b00111111010010101111011010000011;
assign x[  98]= 32'b00111111010001111111011001101010;
assign x[  99]= 32'b00111111010000111111011001010001;
assign x[ 100]= 32'b00111111001111111111011000111001;
assign x[ 101]= 32'b00111111001110111111011000100000;
assign x[ 102]= 32'b00111111001101111111011000000111;
assign x[ 103]= 32'b00111111001100111111010111101110;
assign x[ 104]= 32'b00111111001011111111010111010101;
assign x[ 105]= 32'b00111111001010111111010110111100;
assign x[ 106]= 32'b00111111001001111111010110100100;
assign x[ 107]= 32'b00111111001000111111010110001011;
assign x[ 108]= 32'b00111111000111111111010101110010;
assign x[ 109]= 32'b00111111000110111111010101011001;
assign x[ 110]= 32'b00111111000101111111010101000000;
assign x[ 111]= 32'b00111111000100111111010100101000;
assign x[ 112]= 32'b00111111000011101111010100001111;
assign x[ 113]= 32'b00111111000010101111010011110110;
assign x[ 114]= 32'b00111111000001101111010011011101;
assign x[ 115]= 32'b00111111000000011111010011000101;
assign x[ 116]= 32'b00111110111111011111010010101100;
assign x[ 117]= 32'b00111110111110001111010010010011;
assign x[ 118]= 32'b00111110111101001111010001111011;
assign x[ 119]= 32'b00111110111011111111010001100010;
assign x[ 120]= 32'b00111110111010111111010001001001;
assign x[ 121]= 32'b00111110111001101111010000110000;
assign x[ 122]= 32'b00111110111000011111010000011000;
assign x[ 123]= 32'b00111110110111011111001111111111;
assign x[ 124]= 32'b00111110110110001111001111100110;
assign x[ 125]= 32'b00111110110100111111001111001110;
assign x[ 126]= 32'b00111110110011101111001110110101;
assign x[ 127]= 32'b00111110110010101111001110011100;
assign x[ 128]= 32'b00111110110001011111001110000100;
assign x[ 129]= 32'b00111110110000001111001101101011;
assign x[ 130]= 32'b00111110101110111111001101010010;
assign x[ 131]= 32'b00111110101101101111001100111010;
assign x[ 132]= 32'b00111110101100011111001100100001;
assign x[ 133]= 32'b00111110101011001111001100001000;
assign x[ 134]= 32'b00111110101001111111001011110000;
assign x[ 135]= 32'b00111110101000011111001011010111;
assign x[ 136]= 32'b00111110100111001111001010111111;
assign x[ 137]= 32'b00111110100101111111001010100110;
assign x[ 138]= 32'b00111110100100101111001010001110;
assign x[ 139]= 32'b00111110100011001111001001110101;
assign x[ 140]= 32'b00111110100001111111001001011100;
assign x[ 141]= 32'b00111110100000101111001001000100;
assign x[ 142]= 32'b00111110011111001111001000101011;
assign x[ 143]= 32'b00111110011101111111001000010011;
assign x[ 144]= 32'b00111110011100011111000111111010;
assign x[ 145]= 32'b00111110011011001111000111100010;
assign x[ 146]= 32'b00111110011001101111000111001001;
assign x[ 147]= 32'b00111110011000011111000110110001;
assign x[ 148]= 32'b00111110010110111111000110011000;
assign x[ 149]= 32'b00111110010101011111000110000000;
assign x[ 150]= 32'b00111110010100001111000101100111;
assign x[ 151]= 32'b00111110010010101111000101001111;
assign x[ 152]= 32'b00111110010001001111000100110110;
assign x[ 153]= 32'b00111110001111101111000100011110;
assign x[ 154]= 32'b00111110001110001111000100000101;
assign x[ 155]= 32'b00111110001100111111000011101101;
assign x[ 156]= 32'b00111110001011011111000011010101;
assign x[ 157]= 32'b00111110001001111111000010111100;
assign x[ 158]= 32'b00111110001000011111000010100100;
assign x[ 159]= 32'b00111110000110111111000010001011;
assign x[ 160]= 32'b00111110000101001111000001110011;
assign x[ 161]= 32'b00111110000011101111000001011011;
assign x[ 162]= 32'b00111110000010001111000001000010;
assign x[ 163]= 32'b00111110000000101111000000101010;
assign x[ 164]= 32'b00111101111111001111000000010010;
assign x[ 165]= 32'b00111101111101011110111111111001;
assign x[ 166]= 32'b00111101111011111110111111100001;
assign x[ 167]= 32'b00111101111010011110111111001001;
assign x[ 168]= 32'b00111101111000101110111110110000;
assign x[ 169]= 32'b00111101110111001110111110011000;
assign x[ 170]= 32'b00111101110101101110111110000000;
assign x[ 171]= 32'b00111101110011111110111101100111;
assign x[ 172]= 32'b00111101110010011110111101001111;
assign x[ 173]= 32'b00111101110000101110111100110111;
assign x[ 174]= 32'b00111101101110111110111100011111;
assign x[ 175]= 32'b00111101101101011110111100000110;
assign x[ 176]= 32'b00111101101011101110111011101110;
assign x[ 177]= 32'b00111101101001111110111011010110;
assign x[ 178]= 32'b00111101101000011110111010111110;
assign x[ 179]= 32'b00111101100110101110111010100110;
assign x[ 180]= 32'b00111101100100111110111010001101;
assign x[ 181]= 32'b00111101100011001110111001110101;
assign x[ 182]= 32'b00111101100001011110111001011101;
assign x[ 183]= 32'b00111101011111101110111001000101;
assign x[ 184]= 32'b00111101011101111110111000101101;
assign x[ 185]= 32'b00111101011100001110111000010101;
assign x[ 186]= 32'b00111101011010011110110111111100;
assign x[ 187]= 32'b00111101011000101110110111100100;
assign x[ 188]= 32'b00111101010110111110110111001100;
assign x[ 189]= 32'b00111101010101001110110110110100;
assign x[ 190]= 32'b00111101010011011110110110011100;
assign x[ 191]= 32'b00111101010001011110110110000100;
assign x[ 192]= 32'b00111101001111101110110101101100;
assign x[ 193]= 32'b00111101001101111110110101010100;
assign x[ 194]= 32'b00111101001011111110110100111100;
assign x[ 195]= 32'b00111101001010001110110100100100;
assign x[ 196]= 32'b00111101001000011110110100001100;
assign x[ 197]= 32'b00111101000110011110110011110100;
assign x[ 198]= 32'b00111101000100101110110011011100;
assign x[ 199]= 32'b00111101000010101110110011000100;
assign x[ 200]= 32'b00111101000000101110110010101100;
assign x[ 201]= 32'b00111100111110111110110010010100;
assign x[ 202]= 32'b00111100111100111110110001111100;
assign x[ 203]= 32'b00111100111011001110110001100100;
assign x[ 204]= 32'b00111100111001001110110001001100;
assign x[ 205]= 32'b00111100110111001110110000110100;
assign x[ 206]= 32'b00111100110101001110110000011100;
assign x[ 207]= 32'b00111100110011001110110000000101;
assign x[ 208]= 32'b00111100110001011110101111101101;
assign x[ 209]= 32'b00111100101111011110101111010101;
assign x[ 210]= 32'b00111100101101011110101110111101;
assign x[ 211]= 32'b00111100101011011110101110100101;
assign x[ 212]= 32'b00111100101001011110101110001101;
assign x[ 213]= 32'b00111100100111011110101101110101;
assign x[ 214]= 32'b00111100100101011110101101011110;
assign x[ 215]= 32'b00111100100011001110101101000110;
assign x[ 216]= 32'b00111100100001001110101100101110;
assign x[ 217]= 32'b00111100011111001110101100010110;
assign x[ 218]= 32'b00111100011101001110101011111111;
assign x[ 219]= 32'b00111100011011001110101011100111;
assign x[ 220]= 32'b00111100011000111110101011001111;
assign x[ 221]= 32'b00111100010110111110101010110111;
assign x[ 222]= 32'b00111100010100111110101010100000;
assign x[ 223]= 32'b00111100010010101110101010001000;
assign x[ 224]= 32'b00111100010000101110101001110000;
assign x[ 225]= 32'b00111100001110011110101001011001;
assign x[ 226]= 32'b00111100001100011110101001000001;
assign x[ 227]= 32'b00111100001010001110101000101001;
assign x[ 228]= 32'b00111100001000001110101000010010;
assign x[ 229]= 32'b00111100000101111110100111111010;
assign x[ 230]= 32'b00111100000011101110100111100011;
assign x[ 231]= 32'b00111100000001101110100111001011;
assign x[ 232]= 32'b00111011111111011110100110110100;
assign x[ 233]= 32'b00111011111101001110100110011100;
assign x[ 234]= 32'b00111011111010111110100110000100;
assign x[ 235]= 32'b00111011111000101110100101101101;
assign x[ 236]= 32'b00111011110110101110100101010101;
assign x[ 237]= 32'b00111011110100011110100100111110;
assign x[ 238]= 32'b00111011110010001110100100100110;
assign x[ 239]= 32'b00111011101111111110100100001111;
assign x[ 240]= 32'b00111011101101101110100011110111;
assign x[ 241]= 32'b00111011101011011110100011100000;
assign x[ 242]= 32'b00111011101000111110100011001001;
assign x[ 243]= 32'b00111011100110101110100010110001;
assign x[ 244]= 32'b00111011100100011110100010011010;
assign x[ 245]= 32'b00111011100010001110100010000010;
assign x[ 246]= 32'b00111011011111111110100001101011;
assign x[ 247]= 32'b00111011011101011110100001010100;
assign x[ 248]= 32'b00111011011011001110100000111100;
assign x[ 249]= 32'b00111011011000111110100000100101;
assign x[ 250]= 32'b00111011010110011110100000001110;
assign x[ 251]= 32'b00111011010100001110011111110110;
assign x[ 252]= 32'b00111011010001111110011111011111;
assign x[ 253]= 32'b00111011001111011110011111001000;
assign x[ 254]= 32'b00111011001101001110011110110001;
assign x[ 255]= 32'b00111011001010101110011110011001;
assign x[ 256]= 32'b00111011001000001110011110000010;
assign x[ 257]= 32'b00111011000101111110011101101011;
assign x[ 258]= 32'b00111011000011011110011101010100;
assign x[ 259]= 32'b00111011000000111110011100111101;
assign x[ 260]= 32'b00111010111110101110011100100101;
assign x[ 261]= 32'b00111010111100001110011100001110;
assign x[ 262]= 32'b00111010111001101110011011110111;
assign x[ 263]= 32'b00111010110111001110011011100000;
assign x[ 264]= 32'b00111010110100101110011011001001;
assign x[ 265]= 32'b00111010110010001110011010110010;
assign x[ 266]= 32'b00111010101111101110011010011011;
assign x[ 267]= 32'b00111010101101001110011010000100;
assign x[ 268]= 32'b00111010101010101110011001101101;
assign x[ 269]= 32'b00111010101000001110011001010110;
assign x[ 270]= 32'b00111010100101101110011000111111;
assign x[ 271]= 32'b00111010100011001110011000101000;
assign x[ 272]= 32'b00111010100000101110011000010001;
assign x[ 273]= 32'b00111010011110001110010111111010;
assign x[ 274]= 32'b00111010011011011110010111100011;
assign x[ 275]= 32'b00111010011000111110010111001100;
assign x[ 276]= 32'b00111010010110011110010110110101;
assign x[ 277]= 32'b00111010010011111110010110011110;
assign x[ 278]= 32'b00111010010001001110010110000111;
assign x[ 279]= 32'b00111010001110101110010101110000;
assign x[ 280]= 32'b00111010001011111110010101011001;
assign x[ 281]= 32'b00111010001001011110010101000010;
assign x[ 282]= 32'b00111010000110101110010100101100;
assign x[ 283]= 32'b00111010000100001110010100010101;
assign x[ 284]= 32'b00111010000001011110010011111110;
assign x[ 285]= 32'b00111001111110111110010011100111;
assign x[ 286]= 32'b00111001111100001110010011010000;
assign x[ 287]= 32'b00111001111001011110010010111010;
assign x[ 288]= 32'b00111001110110101110010010100011;
assign x[ 289]= 32'b00111001110100001110010010001100;
assign x[ 290]= 32'b00111001110001011110010001110110;
assign x[ 291]= 32'b00111001101110101110010001011111;
assign x[ 292]= 32'b00111001101011111110010001001000;
assign x[ 293]= 32'b00111001101001001110010000110010;
assign x[ 294]= 32'b00111001100110011110010000011011;
assign x[ 295]= 32'b00111001100011101110010000000100;
assign x[ 296]= 32'b00111001100000111110001111101110;
assign x[ 297]= 32'b00111001011110001110001111010111;
assign x[ 298]= 32'b00111001011011011110001111000001;
assign x[ 299]= 32'b00111001011000101110001110101010;
assign x[ 300]= 32'b00111001010101111110001110010100;
assign x[ 301]= 32'b00111001010011001110001101111101;
assign x[ 302]= 32'b00111001010000011110001101100111;
assign x[ 303]= 32'b00111001001101011110001101010000;
assign x[ 304]= 32'b00111001001010101110001100111010;
assign x[ 305]= 32'b00111001000111111110001100100011;
assign x[ 306]= 32'b00111001000100111110001100001101;
assign x[ 307]= 32'b00111001000010001110001011110110;
assign x[ 308]= 32'b00111000111111011110001011100000;
assign x[ 309]= 32'b00111000111100011110001011001010;
assign x[ 310]= 32'b00111000111001101110001010110011;
assign x[ 311]= 32'b00111000110110101110001010011101;
assign x[ 312]= 32'b00111000110011111110001010000111;
assign x[ 313]= 32'b00111000110000111110001001110000;
assign x[ 314]= 32'b00111000101101111110001001011010;
assign x[ 315]= 32'b00111000101011001110001001000100;
assign x[ 316]= 32'b00111000101000001110001000101101;
assign x[ 317]= 32'b00111000100101001110001000010111;
assign x[ 318]= 32'b00111000100010011110001000000001;
assign x[ 319]= 32'b00111000011111011110000111101011;
assign x[ 320]= 32'b00111000011100011110000111010101;
assign x[ 321]= 32'b00111000011001011110000110111110;
assign x[ 322]= 32'b00111000010110011110000110101000;
assign x[ 323]= 32'b00111000010011011110000110010010;
assign x[ 324]= 32'b00111000010000011110000101111100;
assign x[ 325]= 32'b00111000001101011110000101100110;
assign x[ 326]= 32'b00111000001010011110000101010000;
assign x[ 327]= 32'b00111000000111011110000100111010;
assign x[ 328]= 32'b00111000000100011110000100100100;
assign x[ 329]= 32'b00111000000001011110000100001110;
assign x[ 330]= 32'b00110111111110011110000011111000;
assign x[ 331]= 32'b00110111111011011110000011100010;
assign x[ 332]= 32'b00110111111000001110000011001100;
assign x[ 333]= 32'b00110111110101001110000010110110;
assign x[ 334]= 32'b00110111110010001110000010100000;
assign x[ 335]= 32'b00110111101110111110000010001010;
assign x[ 336]= 32'b00110111101011111110000001110100;
assign x[ 337]= 32'b00110111101000111110000001011110;
assign x[ 338]= 32'b00110111100101101110000001001001;
assign x[ 339]= 32'b00110111100010101110000000110011;
assign x[ 340]= 32'b00110111011111011110000000011101;
assign x[ 341]= 32'b00110111011100011110000000000111;
assign x[ 342]= 32'b00110111011001001101111111110001;
assign x[ 343]= 32'b00110111010101111101111111011100;
assign x[ 344]= 32'b00110111010010111101111111000110;
assign x[ 345]= 32'b00110111001111101101111110110000;
assign x[ 346]= 32'b00110111001100011101111110011011;
assign x[ 347]= 32'b00110111001001011101111110000101;
assign x[ 348]= 32'b00110111000110001101111101101111;
assign x[ 349]= 32'b00110111000010111101111101011010;
assign x[ 350]= 32'b00110110111111101101111101000100;
assign x[ 351]= 32'b00110110111100011101111100101111;
assign x[ 352]= 32'b00110110111001011101111100011001;
assign x[ 353]= 32'b00110110110110001101111100000011;
assign x[ 354]= 32'b00110110110010111101111011101110;
assign x[ 355]= 32'b00110110101111101101111011011000;
assign x[ 356]= 32'b00110110101100011101111011000011;
assign x[ 357]= 32'b00110110101001001101111010101101;
assign x[ 358]= 32'b00110110100101101101111010011000;
assign x[ 359]= 32'b00110110100010011101111010000011;
assign x[ 360]= 32'b00110110011111001101111001101101;
assign x[ 361]= 32'b00110110011011111101111001011000;
assign x[ 362]= 32'b00110110011000101101111001000010;
assign x[ 363]= 32'b00110110010101001101111000101101;
assign x[ 364]= 32'b00110110010001111101111000011000;
assign x[ 365]= 32'b00110110001110101101111000000010;
assign x[ 366]= 32'b00110110001011001101110111101101;
assign x[ 367]= 32'b00110110000111111101110111011000;
assign x[ 368]= 32'b00110110000100101101110111000011;
assign x[ 369]= 32'b00110110000001001101110110101101;
assign x[ 370]= 32'b00110101111101111101110110011000;
assign x[ 371]= 32'b00110101111010011101110110000011;
assign x[ 372]= 32'b00110101110111001101110101101110;
assign x[ 373]= 32'b00110101110011101101110101011001;
assign x[ 374]= 32'b00110101110000001101110101000100;
assign x[ 375]= 32'b00110101101100111101110100101110;
assign x[ 376]= 32'b00110101101001011101110100011001;
assign x[ 377]= 32'b00110101100101111101110100000100;
assign x[ 378]= 32'b00110101100010011101110011101111;
assign x[ 379]= 32'b00110101011111001101110011011010;
assign x[ 380]= 32'b00110101011011101101110011000101;
assign x[ 381]= 32'b00110101011000001101110010110000;
assign x[ 382]= 32'b00110101010100101101110010011011;
assign x[ 383]= 32'b00110101010001001101110010000110;
assign x[ 384]= 32'b00110101001101101101110001110010;
assign x[ 385]= 32'b00110101001010001101110001011101;
assign x[ 386]= 32'b00110101000110101101110001001000;
assign x[ 387]= 32'b00110101000011001101110000110011;
assign x[ 388]= 32'b00110100111111101101110000011110;
assign x[ 389]= 32'b00110100111100001101110000001001;
assign x[ 390]= 32'b00110100111000101101101111110101;
assign x[ 391]= 32'b00110100110101001101101111100000;
assign x[ 392]= 32'b00110100110001101101101111001011;
assign x[ 393]= 32'b00110100101101111101101110110110;
assign x[ 394]= 32'b00110100101010011101101110100010;
assign x[ 395]= 32'b00110100100110111101101110001101;
assign x[ 396]= 32'b00110100100011001101101101111000;
assign x[ 397]= 32'b00110100011111101101101101100100;
assign x[ 398]= 32'b00110100011100001101101101001111;
assign x[ 399]= 32'b00110100011000011101101100111011;
assign x[ 400]= 32'b00110100010100111101101100100110;
assign x[ 401]= 32'b00110100010001001101101100010001;
assign x[ 402]= 32'b00110100001101101101101011111101;
assign x[ 403]= 32'b00110100001001111101101011101000;
assign x[ 404]= 32'b00110100000110011101101011010100;
assign x[ 405]= 32'b00110100000010101101101010111111;
assign x[ 406]= 32'b00110011111110111101101010101011;
assign x[ 407]= 32'b00110011111011011101101010010111;
assign x[ 408]= 32'b00110011110111101101101010000010;
assign x[ 409]= 32'b00110011110011111101101001101110;
assign x[ 410]= 32'b00110011110000011101101001011010;
assign x[ 411]= 32'b00110011101100101101101001000101;
assign x[ 412]= 32'b00110011101000111101101000110001;
assign x[ 413]= 32'b00110011100101001101101000011101;
assign x[ 414]= 32'b00110011100001011101101000001000;
assign x[ 415]= 32'b00110011011101101101100111110100;
assign x[ 416]= 32'b00110011011001111101100111100000;
assign x[ 417]= 32'b00110011010110001101100111001100;
assign x[ 418]= 32'b00110011010010011101100110111000;
assign x[ 419]= 32'b00110011001110101101100110100100;
assign x[ 420]= 32'b00110011001010111101100110001111;
assign x[ 421]= 32'b00110011000111001101100101111011;
assign x[ 422]= 32'b00110011000011011101100101100111;
assign x[ 423]= 32'b00110010111111101101100101010011;
assign x[ 424]= 32'b00110010111011101101100100111111;
assign x[ 425]= 32'b00110010110111111101100100101011;
assign x[ 426]= 32'b00110010110100001101100100010111;
assign x[ 427]= 32'b00110010110000011101100100000011;
assign x[ 428]= 32'b00110010101100011101100011101111;
assign x[ 429]= 32'b00110010101000101101100011011100;
assign x[ 430]= 32'b00110010100100111101100011001000;
assign x[ 431]= 32'b00110010100000111101100010110100;
assign x[ 432]= 32'b00110010011101001101100010100000;
assign x[ 433]= 32'b00110010011001001101100010001100;
assign x[ 434]= 32'b00110010010101011101100001111000;
assign x[ 435]= 32'b00110010010001011101100001100101;
assign x[ 436]= 32'b00110010001101101101100001010001;
assign x[ 437]= 32'b00110010001001101101100000111101;
assign x[ 438]= 32'b00110010000101101101100000101010;
assign x[ 439]= 32'b00110010000001111101100000010110;
assign x[ 440]= 32'b00110001111101111101100000000010;
assign x[ 441]= 32'b00110001111001111101011111101111;
assign x[ 442]= 32'b00110001110110001101011111011011;
assign x[ 443]= 32'b00110001110010001101011111001000;
assign x[ 444]= 32'b00110001101110001101011110110100;
assign x[ 445]= 32'b00110001101010001101011110100000;
assign x[ 446]= 32'b00110001100110001101011110001101;
assign x[ 447]= 32'b00110001100010001101011101111010;
assign x[ 448]= 32'b00110001011110011101011101100110;
assign x[ 449]= 32'b00110001011010011101011101010011;
assign x[ 450]= 32'b00110001010110011101011100111111;
assign x[ 451]= 32'b00110001010010011101011100101100;
assign x[ 452]= 32'b00110001001110001101011100011001;
assign x[ 453]= 32'b00110001001010001101011100000101;
assign x[ 454]= 32'b00110001000110001101011011110010;
assign x[ 455]= 32'b00110001000010001101011011011111;
assign x[ 456]= 32'b00110000111110001101011011001011;
assign x[ 457]= 32'b00110000111010001101011010111000;
assign x[ 458]= 32'b00110000110110001101011010100101;
assign x[ 459]= 32'b00110000110001111101011010010010;
assign x[ 460]= 32'b00110000101101111101011001111111;
assign x[ 461]= 32'b00110000101001111101011001101100;
assign x[ 462]= 32'b00110000100101101101011001011001;
assign x[ 463]= 32'b00110000100001101101011001000101;
assign x[ 464]= 32'b00110000011101101101011000110010;
assign x[ 465]= 32'b00110000011001011101011000011111;
assign x[ 466]= 32'b00110000010101011101011000001100;
assign x[ 467]= 32'b00110000010001001101010111111001;
assign x[ 468]= 32'b00110000001101001101010111100110;
assign x[ 469]= 32'b00110000001000111101010111010100;
assign x[ 470]= 32'b00110000000100111101010111000001;
assign x[ 471]= 32'b00110000000000101101010110101110;
assign x[ 472]= 32'b00101111111100011101010110011011;
assign x[ 473]= 32'b00101111111000011101010110001000;
assign x[ 474]= 32'b00101111110100001101010101110101;
assign x[ 475]= 32'b00101111101111111101010101100011;
assign x[ 476]= 32'b00101111101011111101010101010000;
assign x[ 477]= 32'b00101111100111101101010100111101;
assign x[ 478]= 32'b00101111100011011101010100101010;
assign x[ 479]= 32'b00101111011111001101010100011000;
assign x[ 480]= 32'b00101111011010111101010100000101;
assign x[ 481]= 32'b00101111010110101101010011110011;
assign x[ 482]= 32'b00101111010010011101010011100000;
assign x[ 483]= 32'b00101111001110001101010011001101;
assign x[ 484]= 32'b00101111001010001101010010111011;
assign x[ 485]= 32'b00101111000101101101010010101000;
assign x[ 486]= 32'b00101111000001011101010010010110;
assign x[ 487]= 32'b00101110111101001101010010000011;
assign x[ 488]= 32'b00101110111000111101010001110001;
assign x[ 489]= 32'b00101110110100101101010001011111;
assign x[ 490]= 32'b00101110110000011101010001001100;
assign x[ 491]= 32'b00101110101100001101010000111010;
assign x[ 492]= 32'b00101110100111111101010000101000;
assign x[ 493]= 32'b00101110100011011101010000010101;
assign x[ 494]= 32'b00101110011111001101010000000011;
assign x[ 495]= 32'b00101110011010111101001111110001;
assign x[ 496]= 32'b00101110010110101101001111011111;
assign x[ 497]= 32'b00101110010010001101001111001100;
assign x[ 498]= 32'b00101110001101111101001110111010;
assign x[ 499]= 32'b00101110001001011101001110101000;
assign x[ 500]= 32'b00101110000101001101001110010110;
assign x[ 501]= 32'b00101110000000111101001110000100;
assign x[ 502]= 32'b00101101111100011101001101110010;
assign x[ 503]= 32'b00101101111000001101001101100000;
assign x[ 504]= 32'b00101101110011101101001101001110;
assign x[ 505]= 32'b00101101101111001101001100111100;
assign x[ 506]= 32'b00101101101010111101001100101010;
assign x[ 507]= 32'b00101101100110011101001100011000;
assign x[ 508]= 32'b00101101100010001101001100000110;
assign x[ 509]= 32'b00101101011101101101001011110100;
assign x[ 510]= 32'b00101101011001001101001011100010;
assign x[ 511]= 32'b00101101010100101101001011010001;
assign x[ 512]= 32'b00101101010000011101001010111111;
assign x[ 513]= 32'b00101101001011111101001010101101;
assign x[ 514]= 32'b00101101000111011101001010011011;
assign x[ 515]= 32'b00101101000010111101001010001010;
assign x[ 516]= 32'b00101100111110011101001001111000;
assign x[ 517]= 32'b00101100111010001101001001100110;
assign x[ 518]= 32'b00101100110101101101001001010101;
assign x[ 519]= 32'b00101100110001001101001001000011;
assign x[ 520]= 32'b00101100101100101101001000110001;
assign x[ 521]= 32'b00101100101000001101001000100000;
assign x[ 522]= 32'b00101100100011101101001000001110;
assign x[ 523]= 32'b00101100011111001101000111111101;
assign x[ 524]= 32'b00101100011010101101000111101011;
assign x[ 525]= 32'b00101100010101111101000111011010;
assign x[ 526]= 32'b00101100010001011101000111001001;
assign x[ 527]= 32'b00101100001100111101000110110111;
assign x[ 528]= 32'b00101100001000011101000110100110;
assign x[ 529]= 32'b00101100000011111101000110010101;
assign x[ 530]= 32'b00101011111111001101000110000011;
assign x[ 531]= 32'b00101011111010101101000101110010;
assign x[ 532]= 32'b00101011110110001101000101100001;
assign x[ 533]= 32'b00101011110001101101000101010000;
assign x[ 534]= 32'b00101011101100111101000100111110;
assign x[ 535]= 32'b00101011101000011101000100101101;
assign x[ 536]= 32'b00101011100011101101000100011100;
assign x[ 537]= 32'b00101011011111001101000100001011;
assign x[ 538]= 32'b00101011011010101101000011111010;
assign x[ 539]= 32'b00101011010101111101000011101001;
assign x[ 540]= 32'b00101011010001011101000011011000;
assign x[ 541]= 32'b00101011001100101101000011000111;
assign x[ 542]= 32'b00101011001000001101000010110110;
assign x[ 543]= 32'b00101011000011011101000010100101;
assign x[ 544]= 32'b00101010111110101101000010010100;
assign x[ 545]= 32'b00101010111010001101000010000011;
assign x[ 546]= 32'b00101010110101011101000001110011;
assign x[ 547]= 32'b00101010110000101101000001100010;
assign x[ 548]= 32'b00101010101100001101000001010001;
assign x[ 549]= 32'b00101010100111011101000001000000;
assign x[ 550]= 32'b00101010100010101101000000110000;
assign x[ 551]= 32'b00101010011101111101000000011111;
assign x[ 552]= 32'b00101010011001011101000000001110;
assign x[ 553]= 32'b00101010010100101100111111111110;
assign x[ 554]= 32'b00101010001111111100111111101101;
assign x[ 555]= 32'b00101010001011001100111111011100;
assign x[ 556]= 32'b00101010000110011100111111001100;
assign x[ 557]= 32'b00101010000001101100111110111011;
assign x[ 558]= 32'b00101001111100111100111110101011;
assign x[ 559]= 32'b00101001111000001100111110011010;
assign x[ 560]= 32'b00101001110011011100111110001010;
assign x[ 561]= 32'b00101001101110101100111101111001;
assign x[ 562]= 32'b00101001101001111100111101101001;
assign x[ 563]= 32'b00101001100101001100111101011001;
assign x[ 564]= 32'b00101001100000011100111101001000;
assign x[ 565]= 32'b00101001011011101100111100111000;
assign x[ 566]= 32'b00101001010110101100111100101000;
assign x[ 567]= 32'b00101001010001111100111100011000;
assign x[ 568]= 32'b00101001001101001100111100000111;
assign x[ 569]= 32'b00101001001000011100111011110111;
assign x[ 570]= 32'b00101001000011101100111011100111;
assign x[ 571]= 32'b00101000111110101100111011010111;
assign x[ 572]= 32'b00101000111001111100111011000111;
assign x[ 573]= 32'b00101000110101001100111010110111;
assign x[ 574]= 32'b00101000110000001100111010100111;
assign x[ 575]= 32'b00101000101011011100111010010111;
assign x[ 576]= 32'b00101000100110011100111010000111;
assign x[ 577]= 32'b00101000100001101100111001110111;
assign x[ 578]= 32'b00101000011100101100111001100111;
assign x[ 579]= 32'b00101000010111111100111001010111;
assign x[ 580]= 32'b00101000010010111100111001000111;
assign x[ 581]= 32'b00101000001110001100111000111000;
assign x[ 582]= 32'b00101000001001001100111000101000;
assign x[ 583]= 32'b00101000000100011100111000011000;
assign x[ 584]= 32'b00100111111111011100111000001000;
assign x[ 585]= 32'b00100111111010101100110111111001;
assign x[ 586]= 32'b00100111110101101100110111101001;
assign x[ 587]= 32'b00100111110000101100110111011001;
assign x[ 588]= 32'b00100111101011111100110111001010;
assign x[ 589]= 32'b00100111100110111100110110111010;
assign x[ 590]= 32'b00100111100001111100110110101011;
assign x[ 591]= 32'b00100111011100111100110110011011;
assign x[ 592]= 32'b00100111010111111100110110001100;
assign x[ 593]= 32'b00100111010011001100110101111100;
assign x[ 594]= 32'b00100111001110001100110101101101;
assign x[ 595]= 32'b00100111001001001100110101011101;
assign x[ 596]= 32'b00100111000100001100110101001110;
assign x[ 597]= 32'b00100110111111001100110100111111;
assign x[ 598]= 32'b00100110111010001100110100110000;
assign x[ 599]= 32'b00100110110101001100110100100000;
assign x[ 600]= 32'b00100110110000001100110100010001;
assign x[ 601]= 32'b00100110101011001100110100000010;
assign x[ 602]= 32'b00100110100110001100110011110011;
assign x[ 603]= 32'b00100110100001001100110011100011;
assign x[ 604]= 32'b00100110011100001100110011010100;
assign x[ 605]= 32'b00100110010111001100110011000101;
assign x[ 606]= 32'b00100110010010001100110010110110;
assign x[ 607]= 32'b00100110001101001100110010100111;
assign x[ 608]= 32'b00100110000111111100110010011000;
assign x[ 609]= 32'b00100110000010111100110010001001;
assign x[ 610]= 32'b00100101111101111100110001111010;
assign x[ 611]= 32'b00100101111000111100110001101011;
assign x[ 612]= 32'b00100101110011111100110001011101;
assign x[ 613]= 32'b00100101101110101100110001001110;
assign x[ 614]= 32'b00100101101001101100110000111111;
assign x[ 615]= 32'b00100101100100101100110000110000;
assign x[ 616]= 32'b00100101011111011100110000100001;
assign x[ 617]= 32'b00100101011010011100110000010011;
assign x[ 618]= 32'b00100101010101001100110000000100;
assign x[ 619]= 32'b00100101010000001100101111110101;
assign x[ 620]= 32'b00100101001011001100101111100111;
assign x[ 621]= 32'b00100101000101111100101111011000;
assign x[ 622]= 32'b00100101000000111100101111001010;
assign x[ 623]= 32'b00100100111011101100101110111011;
assign x[ 624]= 32'b00100100110110101100101110101101;
assign x[ 625]= 32'b00100100110001011100101110011110;
assign x[ 626]= 32'b00100100101100001100101110010000;
assign x[ 627]= 32'b00100100100111001100101110000001;
assign x[ 628]= 32'b00100100100001111100101101110011;
assign x[ 629]= 32'b00100100011100111100101101100101;
assign x[ 630]= 32'b00100100010111101100101101010110;
assign x[ 631]= 32'b00100100010010011100101101001000;
assign x[ 632]= 32'b00100100001101001100101100111010;
assign x[ 633]= 32'b00100100001000001100101100101100;
assign x[ 634]= 32'b00100100000010111100101100011110;
assign x[ 635]= 32'b00100011111101101100101100001111;
assign x[ 636]= 32'b00100011111000011100101100000001;
assign x[ 637]= 32'b00100011110011011100101011110011;
assign x[ 638]= 32'b00100011101110001100101011100101;
assign x[ 639]= 32'b00100011101000111100101011010111;
assign x[ 640]= 32'b00100011100011101100101011001001;
assign x[ 641]= 32'b00100011011110011100101010111011;
assign x[ 642]= 32'b00100011011001001100101010101101;
assign x[ 643]= 32'b00100011010011111100101010011111;
assign x[ 644]= 32'b00100011001110101100101010010010;
assign x[ 645]= 32'b00100011001001011100101010000100;
assign x[ 646]= 32'b00100011000100001100101001110110;
assign x[ 647]= 32'b00100010111110111100101001101000;
assign x[ 648]= 32'b00100010111001101100101001011011;
assign x[ 649]= 32'b00100010110100011100101001001101;
assign x[ 650]= 32'b00100010101111001100101000111111;
assign x[ 651]= 32'b00100010101001111100101000110010;
assign x[ 652]= 32'b00100010100100101100101000100100;
assign x[ 653]= 32'b00100010011111011100101000010110;
assign x[ 654]= 32'b00100010011001111100101000001001;
assign x[ 655]= 32'b00100010010100101100100111111011;
assign x[ 656]= 32'b00100010001111011100100111101110;
assign x[ 657]= 32'b00100010001010001100100111100000;
assign x[ 658]= 32'b00100010000100101100100111010011;
assign x[ 659]= 32'b00100001111111011100100111000110;
assign x[ 660]= 32'b00100001111010001100100110111000;
assign x[ 661]= 32'b00100001110100101100100110101011;
assign x[ 662]= 32'b00100001101111011100100110011110;
assign x[ 663]= 32'b00100001101010001100100110010001;
assign x[ 664]= 32'b00100001100100101100100110000011;
assign x[ 665]= 32'b00100001011111011100100101110110;
assign x[ 666]= 32'b00100001011010001100100101101001;
assign x[ 667]= 32'b00100001010100101100100101011100;
assign x[ 668]= 32'b00100001001111011100100101001111;
assign x[ 669]= 32'b00100001001001111100100101000010;
assign x[ 670]= 32'b00100001000100101100100100110101;
assign x[ 671]= 32'b00100000111111001100100100101000;
assign x[ 672]= 32'b00100000111001111100100100011011;
assign x[ 673]= 32'b00100000110100011100100100001110;
assign x[ 674]= 32'b00100000101110111100100100000001;
assign x[ 675]= 32'b00100000101001101100100011110100;
assign x[ 676]= 32'b00100000100100001100100011101000;
assign x[ 677]= 32'b00100000011110111100100011011011;
assign x[ 678]= 32'b00100000011001011100100011001110;
assign x[ 679]= 32'b00100000010011111100100011000001;
assign x[ 680]= 32'b00100000001110011100100010110101;
assign x[ 681]= 32'b00100000001001001100100010101000;
assign x[ 682]= 32'b00100000000011101100100010011011;
assign x[ 683]= 32'b00011111111110001100100010001111;
assign x[ 684]= 32'b00011111111000101100100010000010;
assign x[ 685]= 32'b00011111110011011100100001110110;
assign x[ 686]= 32'b00011111101101111100100001101001;
assign x[ 687]= 32'b00011111101000011100100001011101;
assign x[ 688]= 32'b00011111100010111100100001010000;
assign x[ 689]= 32'b00011111011101011100100001000100;
assign x[ 690]= 32'b00011111010111111100100000111000;
assign x[ 691]= 32'b00011111010010011100100000101011;
assign x[ 692]= 32'b00011111001101001100100000011111;
assign x[ 693]= 32'b00011111000111101100100000010011;
assign x[ 694]= 32'b00011111000010001100100000000111;
assign x[ 695]= 32'b00011110111100101100011111111011;
assign x[ 696]= 32'b00011110110111001100011111101110;
assign x[ 697]= 32'b00011110110001101100011111100010;
assign x[ 698]= 32'b00011110101100001100011111010110;
assign x[ 699]= 32'b00011110100110011100011111001010;
assign x[ 700]= 32'b00011110100000111100011110111110;
assign x[ 701]= 32'b00011110011011011100011110110010;
assign x[ 702]= 32'b00011110010101111100011110100110;
assign x[ 703]= 32'b00011110010000011100011110011010;
assign x[ 704]= 32'b00011110001010111100011110001111;
assign x[ 705]= 32'b00011110000101011100011110000011;
assign x[ 706]= 32'b00011101111111101100011101110111;
assign x[ 707]= 32'b00011101111010001100011101101011;
assign x[ 708]= 32'b00011101110100101100011101011111;
assign x[ 709]= 32'b00011101101111001100011101010100;
assign x[ 710]= 32'b00011101101001101100011101001000;
assign x[ 711]= 32'b00011101100011111100011100111101;
assign x[ 712]= 32'b00011101011110011100011100110001;
assign x[ 713]= 32'b00011101011000111100011100100101;
assign x[ 714]= 32'b00011101010011001100011100011010;
assign x[ 715]= 32'b00011101001101101100011100001110;
assign x[ 716]= 32'b00011101001000001100011100000011;
assign x[ 717]= 32'b00011101000010011100011011110111;
assign x[ 718]= 32'b00011100111100111100011011101100;
assign x[ 719]= 32'b00011100110111001100011011100001;
assign x[ 720]= 32'b00011100110001101100011011010101;
assign x[ 721]= 32'b00011100101011111100011011001010;
assign x[ 722]= 32'b00011100100110011100011010111111;
assign x[ 723]= 32'b00011100100000111100011010110100;
assign x[ 724]= 32'b00011100011011001100011010101000;
assign x[ 725]= 32'b00011100010101011100011010011101;
assign x[ 726]= 32'b00011100001111111100011010010010;
assign x[ 727]= 32'b00011100001010001100011010000111;
assign x[ 728]= 32'b00011100000100101100011001111100;
assign x[ 729]= 32'b00011011111110111100011001110001;
assign x[ 730]= 32'b00011011111001011100011001100110;
assign x[ 731]= 32'b00011011110011101100011001011011;
assign x[ 732]= 32'b00011011101101111100011001010000;
assign x[ 733]= 32'b00011011101000011100011001000101;
assign x[ 734]= 32'b00011011100010101100011000111011;
assign x[ 735]= 32'b00011011011100111100011000110000;
assign x[ 736]= 32'b00011011010111011100011000100101;
assign x[ 737]= 32'b00011011010001101100011000011010;
assign x[ 738]= 32'b00011011001011111100011000010000;
assign x[ 739]= 32'b00011011000110001100011000000101;
assign x[ 740]= 32'b00011011000000101100010111111010;
assign x[ 741]= 32'b00011010111010111100010111110000;
assign x[ 742]= 32'b00011010110101001100010111100101;
assign x[ 743]= 32'b00011010101111011100010111011011;
assign x[ 744]= 32'b00011010101001101100010111010000;
assign x[ 745]= 32'b00011010100011111100010111000110;
assign x[ 746]= 32'b00011010011110011100010110111011;
assign x[ 747]= 32'b00011010011000101100010110110001;
assign x[ 748]= 32'b00011010010010111100010110100111;
assign x[ 749]= 32'b00011010001101001100010110011100;
assign x[ 750]= 32'b00011010000111011100010110010010;
assign x[ 751]= 32'b00011010000001101100010110001000;
assign x[ 752]= 32'b00011001111011111100010101111110;
assign x[ 753]= 32'b00011001110110001100010101110011;
assign x[ 754]= 32'b00011001110000011100010101101001;
assign x[ 755]= 32'b00011001101010101100010101011111;
assign x[ 756]= 32'b00011001100100111100010101010101;
assign x[ 757]= 32'b00011001011111001100010101001011;
assign x[ 758]= 32'b00011001011001011100010101000001;
assign x[ 759]= 32'b00011001010011101100010100110111;
assign x[ 760]= 32'b00011001001101111100010100101101;
assign x[ 761]= 32'b00011001001000001100010100100011;
assign x[ 762]= 32'b00011001000010001100010100011010;
assign x[ 763]= 32'b00011000111100011100010100010000;
assign x[ 764]= 32'b00011000110110101100010100000110;
assign x[ 765]= 32'b00011000110000111100010011111100;
assign x[ 766]= 32'b00011000101011001100010011110010;
assign x[ 767]= 32'b00011000100101011100010011101001;
assign x[ 768]= 32'b00011000011111011100010011011111;
assign x[ 769]= 32'b00011000011001101100010011010110;
assign x[ 770]= 32'b00011000010011111100010011001100;
assign x[ 771]= 32'b00011000001110001100010011000010;
assign x[ 772]= 32'b00011000001000001100010010111001;
assign x[ 773]= 32'b00011000000010011100010010110000;
assign x[ 774]= 32'b00010111111100101100010010100110;
assign x[ 775]= 32'b00010111110110101100010010011101;
assign x[ 776]= 32'b00010111110000111100010010010011;
assign x[ 777]= 32'b00010111101011001100010010001010;
assign x[ 778]= 32'b00010111100101001100010010000001;
assign x[ 779]= 32'b00010111011111011100010001111000;
assign x[ 780]= 32'b00010111011001101100010001101110;
assign x[ 781]= 32'b00010111010011101100010001100101;
assign x[ 782]= 32'b00010111001101111100010001011100;
assign x[ 783]= 32'b00010111000111111100010001010011;
assign x[ 784]= 32'b00010111000010001100010001001010;
assign x[ 785]= 32'b00010110111100011100010001000001;
assign x[ 786]= 32'b00010110110110011100010000111000;
assign x[ 787]= 32'b00010110110000101100010000101111;
assign x[ 788]= 32'b00010110101010101100010000100110;
assign x[ 789]= 32'b00010110100100111100010000011101;
assign x[ 790]= 32'b00010110011110111100010000010100;
assign x[ 791]= 32'b00010110011001001100010000001011;
assign x[ 792]= 32'b00010110010011001100010000000011;
assign x[ 793]= 32'b00010110001101001100001111111010;
assign x[ 794]= 32'b00010110000111011100001111110001;
assign x[ 795]= 32'b00010110000001011100001111101001;
assign x[ 796]= 32'b00010101111011101100001111100000;
assign x[ 797]= 32'b00010101110101101100001111010111;
assign x[ 798]= 32'b00010101101111101100001111001111;
assign x[ 799]= 32'b00010101101001111100001111000110;
assign x[ 800]= 32'b00010101100011111100001110111110;
assign x[ 801]= 32'b00010101011101111100001110110101;
assign x[ 802]= 32'b00010101011000001100001110101101;
assign x[ 803]= 32'b00010101010010001100001110100101;
assign x[ 804]= 32'b00010101001100001100001110011100;
assign x[ 805]= 32'b00010101000110011100001110010100;
assign x[ 806]= 32'b00010101000000011100001110001100;
assign x[ 807]= 32'b00010100111010011100001110000011;
assign x[ 808]= 32'b00010100110100011100001101111011;
assign x[ 809]= 32'b00010100101110101100001101110011;
assign x[ 810]= 32'b00010100101000101100001101101011;
assign x[ 811]= 32'b00010100100010101100001101100011;
assign x[ 812]= 32'b00010100011100101100001101011011;
assign x[ 813]= 32'b00010100010110101100001101010011;
assign x[ 814]= 32'b00010100010000111100001101001011;
assign x[ 815]= 32'b00010100001010111100001101000011;
assign x[ 816]= 32'b00010100000100111100001100111011;
assign x[ 817]= 32'b00010011111110111100001100110011;
assign x[ 818]= 32'b00010011111000111100001100101011;
assign x[ 819]= 32'b00010011110010111100001100100011;
assign x[ 820]= 32'b00010011101100111100001100011100;
assign x[ 821]= 32'b00010011100110111100001100010100;
assign x[ 822]= 32'b00010011100000111100001100001100;
assign x[ 823]= 32'b00010011011011001100001100000101;
assign x[ 824]= 32'b00010011010101001100001011111101;
assign x[ 825]= 32'b00010011001111001100001011110101;
assign x[ 826]= 32'b00010011001001001100001011101110;
assign x[ 827]= 32'b00010011000011001100001011100110;
assign x[ 828]= 32'b00010010111101001100001011011111;
assign x[ 829]= 32'b00010010110111001100001011011000;
assign x[ 830]= 32'b00010010110001001100001011010000;
assign x[ 831]= 32'b00010010101011001100001011001001;
assign x[ 832]= 32'b00010010100101001100001011000001;
assign x[ 833]= 32'b00010010011110111100001010111010;
assign x[ 834]= 32'b00010010011000111100001010110011;
assign x[ 835]= 32'b00010010010010111100001010101100;
assign x[ 836]= 32'b00010010001100111100001010100101;
assign x[ 837]= 32'b00010010000110111100001010011101;
assign x[ 838]= 32'b00010010000000111100001010010110;
assign x[ 839]= 32'b00010001111010111100001010001111;
assign x[ 840]= 32'b00010001110100111100001010001000;
assign x[ 841]= 32'b00010001101110111100001010000001;
assign x[ 842]= 32'b00010001101000101100001001111010;
assign x[ 843]= 32'b00010001100010101100001001110011;
assign x[ 844]= 32'b00010001011100101100001001101101;
assign x[ 845]= 32'b00010001010110101100001001100110;
assign x[ 846]= 32'b00010001010000101100001001011111;
assign x[ 847]= 32'b00010001001010101100001001011000;
assign x[ 848]= 32'b00010001000100011100001001010001;
assign x[ 849]= 32'b00010000111110011100001001001011;
assign x[ 850]= 32'b00010000111000011100001001000100;
assign x[ 851]= 32'b00010000110010011100001000111110;
assign x[ 852]= 32'b00010000101100001100001000110111;
assign x[ 853]= 32'b00010000100110001100001000110000;
assign x[ 854]= 32'b00010000100000001100001000101010;
assign x[ 855]= 32'b00010000011010001100001000100011;
assign x[ 856]= 32'b00010000010011111100001000011101;
assign x[ 857]= 32'b00010000001101111100001000010111;
assign x[ 858]= 32'b00010000000111111100001000010000;
assign x[ 859]= 32'b00010000000001101100001000001010;
assign x[ 860]= 32'b00001111111011101100001000000100;
assign x[ 861]= 32'b00001111110101101100000111111101;
assign x[ 862]= 32'b00001111101111011100000111110111;
assign x[ 863]= 32'b00001111101001011100000111110001;
assign x[ 864]= 32'b00001111100011001100000111101011;
assign x[ 865]= 32'b00001111011101001100000111100101;
assign x[ 866]= 32'b00001111010111001100000111011111;
assign x[ 867]= 32'b00001111010000111100000111011001;
assign x[ 868]= 32'b00001111001010111100000111010011;
assign x[ 869]= 32'b00001111000100101100000111001101;
assign x[ 870]= 32'b00001110111110101100000111000111;
assign x[ 871]= 32'b00001110111000101100000111000001;
assign x[ 872]= 32'b00001110110010011100000110111011;
assign x[ 873]= 32'b00001110101100011100000110110110;
assign x[ 874]= 32'b00001110100110001100000110110000;
assign x[ 875]= 32'b00001110100000001100000110101010;
assign x[ 876]= 32'b00001110011001111100000110100100;
assign x[ 877]= 32'b00001110010011111100000110011111;
assign x[ 878]= 32'b00001110001101101100000110011001;
assign x[ 879]= 32'b00001110000111101100000110010100;
assign x[ 880]= 32'b00001110000001011100000110001110;
assign x[ 881]= 32'b00001101111011011100000110001001;
assign x[ 882]= 32'b00001101110101001100000110000011;
assign x[ 883]= 32'b00001101101111001100000101111110;
assign x[ 884]= 32'b00001101101000111100000101111000;
assign x[ 885]= 32'b00001101100010111100000101110011;
assign x[ 886]= 32'b00001101011100101100000101101110;
assign x[ 887]= 32'b00001101010110011100000101101000;
assign x[ 888]= 32'b00001101010000011100000101100011;
assign x[ 889]= 32'b00001101001010001100000101011110;
assign x[ 890]= 32'b00001101000100001100000101011001;
assign x[ 891]= 32'b00001100111101111100000101010100;
assign x[ 892]= 32'b00001100110111101100000101001111;
assign x[ 893]= 32'b00001100110001101100000101001010;
assign x[ 894]= 32'b00001100101011011100000101000101;
assign x[ 895]= 32'b00001100100101011100000101000000;
assign x[ 896]= 32'b00001100011111001100000100111011;
assign x[ 897]= 32'b00001100011000111100000100110110;
assign x[ 898]= 32'b00001100010010111100000100110001;
assign x[ 899]= 32'b00001100001100101100000100101100;
assign x[ 900]= 32'b00001100000110011100000100101000;
assign x[ 901]= 32'b00001100000000011100000100100011;
assign x[ 902]= 32'b00001011111010001100000100011110;
assign x[ 903]= 32'b00001011110011111100000100011001;
assign x[ 904]= 32'b00001011101101101100000100010101;
assign x[ 905]= 32'b00001011100111101100000100010000;
assign x[ 906]= 32'b00001011100001011100000100001100;
assign x[ 907]= 32'b00001011011011001100000100000111;
assign x[ 908]= 32'b00001011010101001100000100000011;
assign x[ 909]= 32'b00001011001110111100000011111110;
assign x[ 910]= 32'b00001011001000101100000011111010;
assign x[ 911]= 32'b00001011000010011100000011110110;
assign x[ 912]= 32'b00001010111100011100000011110001;
assign x[ 913]= 32'b00001010110110001100000011101101;
assign x[ 914]= 32'b00001010101111111100000011101001;
assign x[ 915]= 32'b00001010101001101100000011100100;
assign x[ 916]= 32'b00001010100011011100000011100000;
assign x[ 917]= 32'b00001010011101011100000011011100;
assign x[ 918]= 32'b00001010010111001100000011011000;
assign x[ 919]= 32'b00001010010000111100000011010100;
assign x[ 920]= 32'b00001010001010101100000011010000;
assign x[ 921]= 32'b00001010000100011100000011001100;
assign x[ 922]= 32'b00001001111110011100000011001000;
assign x[ 923]= 32'b00001001111000001100000011000100;
assign x[ 924]= 32'b00001001110001111100000011000000;
assign x[ 925]= 32'b00001001101011101100000010111101;
assign x[ 926]= 32'b00001001100101011100000010111001;
assign x[ 927]= 32'b00001001011111001100000010110101;
assign x[ 928]= 32'b00001001011001001100000010110001;
assign x[ 929]= 32'b00001001010010111100000010101110;
assign x[ 930]= 32'b00001001001100101100000010101010;
assign x[ 931]= 32'b00001001000110011100000010100110;
assign x[ 932]= 32'b00001001000000001100000010100011;
assign x[ 933]= 32'b00001000111001111100000010011111;
assign x[ 934]= 32'b00001000110011101100000010011100;
assign x[ 935]= 32'b00001000101101011100000010011000;
assign x[ 936]= 32'b00001000100111001100000010010101;
assign x[ 937]= 32'b00001000100001001100000010010010;
assign x[ 938]= 32'b00001000011010111100000010001110;
assign x[ 939]= 32'b00001000010100101100000010001011;
assign x[ 940]= 32'b00001000001110011100000010001000;
assign x[ 941]= 32'b00001000001000001100000010000101;
assign x[ 942]= 32'b00001000000001111100000010000001;
assign x[ 943]= 32'b00000111111011101100000001111110;
assign x[ 944]= 32'b00000111110101011100000001111011;
assign x[ 945]= 32'b00000111101111001100000001111000;
assign x[ 946]= 32'b00000111101000111100000001110101;
assign x[ 947]= 32'b00000111100010101100000001110010;
assign x[ 948]= 32'b00000111011100011100000001101111;
assign x[ 949]= 32'b00000111010110001100000001101100;
assign x[ 950]= 32'b00000111001111111100000001101001;
assign x[ 951]= 32'b00000111001001101100000001100111;
assign x[ 952]= 32'b00000111000011011100000001100100;
assign x[ 953]= 32'b00000110111101001100000001100001;
assign x[ 954]= 32'b00000110110110111100000001011110;
assign x[ 955]= 32'b00000110110000101100000001011100;
assign x[ 956]= 32'b00000110101010011100000001011001;
assign x[ 957]= 32'b00000110100100001100000001010110;
assign x[ 958]= 32'b00000110011101111100000001010100;
assign x[ 959]= 32'b00000110010111101100000001010001;
assign x[ 960]= 32'b00000110010001011100000001001111;
assign x[ 961]= 32'b00000110001011001100000001001100;
assign x[ 962]= 32'b00000110000100111100000001001010;
assign x[ 963]= 32'b00000101111110101100000001001000;
assign x[ 964]= 32'b00000101111000011100000001000101;
assign x[ 965]= 32'b00000101110010001100000001000011;
assign x[ 966]= 32'b00000101101011111100000001000001;
assign x[ 967]= 32'b00000101100101101100000000111111;
assign x[ 968]= 32'b00000101011111011100000000111100;
assign x[ 969]= 32'b00000101011001001100000000111010;
assign x[ 970]= 32'b00000101010010111100000000111000;
assign x[ 971]= 32'b00000101001100101100000000110110;
assign x[ 972]= 32'b00000101000110011100000000110100;
assign x[ 973]= 32'b00000101000000001100000000110010;
assign x[ 974]= 32'b00000100111001111100000000110000;
assign x[ 975]= 32'b00000100110011101100000000101110;
assign x[ 976]= 32'b00000100101101011100000000101100;
assign x[ 977]= 32'b00000100100111001100000000101011;
assign x[ 978]= 32'b00000100100000111100000000101001;
assign x[ 979]= 32'b00000100011010101100000000100111;
assign x[ 980]= 32'b00000100010100011100000000100101;
assign x[ 981]= 32'b00000100001101111100000000100100;
assign x[ 982]= 32'b00000100000111101100000000100010;
assign x[ 983]= 32'b00000100000001011100000000100000;
assign x[ 984]= 32'b00000011111011001100000000011111;
assign x[ 985]= 32'b00000011110100111100000000011101;
assign x[ 986]= 32'b00000011101110101100000000011100;
assign x[ 987]= 32'b00000011101000011100000000011010;
assign x[ 988]= 32'b00000011100010001100000000011001;
assign x[ 989]= 32'b00000011011011111100000000011000;
assign x[ 990]= 32'b00000011010101101100000000010110;
assign x[ 991]= 32'b00000011001111011100000000010101;
assign x[ 992]= 32'b00000011001000111100000000010100;
assign x[ 993]= 32'b00000011000010101100000000010011;
assign x[ 994]= 32'b00000010111100011100000000010001;
assign x[ 995]= 32'b00000010110110001100000000010000;
assign x[ 996]= 32'b00000010101111111100000000001111;
assign x[ 997]= 32'b00000010101001101100000000001110;
assign x[ 998]= 32'b00000010100011011100000000001101;
assign x[ 999]= 32'b00000010011101001100000000001100;
assign x[1000]= 32'b00000010010110111100000000001011;
assign x[1001]= 32'b00000010010000011100000000001010;
assign x[1002]= 32'b00000010001010001100000000001001;
assign x[1003]= 32'b00000010000011111100000000001001;
assign x[1004]= 32'b00000001111101101100000000001000;
assign x[1005]= 32'b00000001110111011100000000000111;
assign x[1006]= 32'b00000001110001001100000000000110;
assign x[1007]= 32'b00000001101010111100000000000110;
assign x[1008]= 32'b00000001100100101100000000000101;
assign x[1009]= 32'b00000001011110001100000000000100;
assign x[1010]= 32'b00000001010111111100000000000100;
assign x[1011]= 32'b00000001010001101100000000000011;
assign x[1012]= 32'b00000001001011011100000000000011;
assign x[1013]= 32'b00000001000101001100000000000010;
assign x[1014]= 32'b00000000111110111100000000000010;
assign x[1015]= 32'b00000000111000101100000000000010;
assign x[1016]= 32'b00000000110010011100000000000001;
assign x[1017]= 32'b00000000101011111100000000000001;
assign x[1018]= 32'b00000000100101101100000000000001;
assign x[1019]= 32'b00000000011111011100000000000000;
assign x[1020]= 32'b00000000011001001100000000000000;
assign x[1021]= 32'b00000000010010111100000000000000;
assign x[1022]= 32'b00000000001100101100000000000000;
assign x[1023]= 32'b00000000000110011100000000000000;
assign x[1024]= 32'b00000000000000001100000000000000;
assign x[1025]= 32'b11111111111001111100000000000000;
assign x[1026]= 32'b11111111110011101100000000000000;
assign x[1027]= 32'b11111111101101011100000000000000;
assign x[1028]= 32'b11111111100110111100000000000000;
assign x[1029]= 32'b11111111100000101100000000000000;
assign x[1030]= 32'b11111111011010011100000000000001;
assign x[1031]= 32'b11111111010100001100000000000001;
assign x[1032]= 32'b11111111001101111100000000000001;
assign x[1033]= 32'b11111111000111101100000000000010;
assign x[1034]= 32'b11111111000001011100000000000010;
assign x[1035]= 32'b11111110111011001100000000000010;
assign x[1036]= 32'b11111110110100101100000000000011;
assign x[1037]= 32'b11111110101110011100000000000011;
assign x[1038]= 32'b11111110101000001100000000000100;
assign x[1039]= 32'b11111110100001111100000000000100;
assign x[1040]= 32'b11111110011011101100000000000101;
assign x[1041]= 32'b11111110010101011100000000000110;
assign x[1042]= 32'b11111110001111001100000000000110;
assign x[1043]= 32'b11111110001000111100000000000111;
assign x[1044]= 32'b11111110000010011100000000001000;
assign x[1045]= 32'b11111101111100001100000000001001;
assign x[1046]= 32'b11111101110101111100000000001001;
assign x[1047]= 32'b11111101101111101100000000001010;
assign x[1048]= 32'b11111101101001011100000000001011;
assign x[1049]= 32'b11111101100011001100000000001100;
assign x[1050]= 32'b11111101011100111100000000001101;
assign x[1051]= 32'b11111101010110101100000000001110;
assign x[1052]= 32'b11111101010000001100000000001111;
assign x[1053]= 32'b11111101001001111100000000010000;
assign x[1054]= 32'b11111101000011101100000000010001;
assign x[1055]= 32'b11111100111101011100000000010011;
assign x[1056]= 32'b11111100110111001100000000010100;
assign x[1057]= 32'b11111100110000111100000000010101;
assign x[1058]= 32'b11111100101010101100000000010110;
assign x[1059]= 32'b11111100100100011100000000011000;
assign x[1060]= 32'b11111100011110001100000000011001;
assign x[1061]= 32'b11111100010111111100000000011010;
assign x[1062]= 32'b11111100010001011100000000011100;
assign x[1063]= 32'b11111100001011001100000000011101;
assign x[1064]= 32'b11111100000100111100000000011111;
assign x[1065]= 32'b11111011111110101100000000100000;
assign x[1066]= 32'b11111011111000011100000000100010;
assign x[1067]= 32'b11111011110010001100000000100100;
assign x[1068]= 32'b11111011101011111100000000100101;
assign x[1069]= 32'b11111011100101101100000000100111;
assign x[1070]= 32'b11111011011111011100000000101001;
assign x[1071]= 32'b11111011011001001100000000101011;
assign x[1072]= 32'b11111011010010111100000000101100;
assign x[1073]= 32'b11111011001100101100000000101110;
assign x[1074]= 32'b11111011000110011100000000110000;
assign x[1075]= 32'b11111011000000001100000000110010;
assign x[1076]= 32'b11111010111001101100000000110100;
assign x[1077]= 32'b11111010110011011100000000110110;
assign x[1078]= 32'b11111010101101001100000000111000;
assign x[1079]= 32'b11111010100110111100000000111010;
assign x[1080]= 32'b11111010100000101100000000111100;
assign x[1081]= 32'b11111010011010011100000000111111;
assign x[1082]= 32'b11111010010100001100000001000001;
assign x[1083]= 32'b11111010001101111100000001000011;
assign x[1084]= 32'b11111010000111101100000001000101;
assign x[1085]= 32'b11111010000001011100000001001000;
assign x[1086]= 32'b11111001111011001100000001001010;
assign x[1087]= 32'b11111001110100111100000001001100;
assign x[1088]= 32'b11111001101110101100000001001111;
assign x[1089]= 32'b11111001101000011100000001010001;
assign x[1090]= 32'b11111001100010001100000001010100;
assign x[1091]= 32'b11111001011011111100000001010110;
assign x[1092]= 32'b11111001010101101100000001011001;
assign x[1093]= 32'b11111001001111011100000001011100;
assign x[1094]= 32'b11111001001001001100000001011110;
assign x[1095]= 32'b11111001000010111100000001100001;
assign x[1096]= 32'b11111000111100101100000001100100;
assign x[1097]= 32'b11111000110110011100000001100111;
assign x[1098]= 32'b11111000110000001100000001101001;
assign x[1099]= 32'b11111000101001111100000001101100;
assign x[1100]= 32'b11111000100011101100000001101111;
assign x[1101]= 32'b11111000011101011100000001110010;
assign x[1102]= 32'b11111000010111001100000001110101;
assign x[1103]= 32'b11111000010000111100000001111000;
assign x[1104]= 32'b11111000001010101100000001111011;
assign x[1105]= 32'b11111000000100011100000001111110;
assign x[1106]= 32'b11110111111110011100000010000001;
assign x[1107]= 32'b11110111111000001100000010000101;
assign x[1108]= 32'b11110111110001111100000010001000;
assign x[1109]= 32'b11110111101011101100000010001011;
assign x[1110]= 32'b11110111100101011100000010001110;
assign x[1111]= 32'b11110111011111001100000010010010;
assign x[1112]= 32'b11110111011000111100000010010101;
assign x[1113]= 32'b11110111010010101100000010011000;
assign x[1114]= 32'b11110111001100011100000010011100;
assign x[1115]= 32'b11110111000110001100000010011111;
assign x[1116]= 32'b11110110111111111100000010100011;
assign x[1117]= 32'b11110110111001111100000010100110;
assign x[1118]= 32'b11110110110011101100000010101010;
assign x[1119]= 32'b11110110101101011100000010101110;
assign x[1120]= 32'b11110110100111001100000010110001;
assign x[1121]= 32'b11110110100000111100000010110101;
assign x[1122]= 32'b11110110011010101100000010111001;
assign x[1123]= 32'b11110110010100011100000010111101;
assign x[1124]= 32'b11110110001110011100000011000000;
assign x[1125]= 32'b11110110001000001100000011000100;
assign x[1126]= 32'b11110110000001111100000011001000;
assign x[1127]= 32'b11110101111011101100000011001100;
assign x[1128]= 32'b11110101110101011100000011010000;
assign x[1129]= 32'b11110101101111001100000011010100;
assign x[1130]= 32'b11110101101001001100000011011000;
assign x[1131]= 32'b11110101100010111100000011011100;
assign x[1132]= 32'b11110101011100101100000011100000;
assign x[1133]= 32'b11110101010110011100000011100100;
assign x[1134]= 32'b11110101010000001100000011101001;
assign x[1135]= 32'b11110101001010001100000011101101;
assign x[1136]= 32'b11110101000011111100000011110001;
assign x[1137]= 32'b11110100111101101100000011110110;
assign x[1138]= 32'b11110100110111011100000011111010;
assign x[1139]= 32'b11110100110001011100000011111110;
assign x[1140]= 32'b11110100101011001100000100000011;
assign x[1141]= 32'b11110100100100111100000100000111;
assign x[1142]= 32'b11110100011110111100000100001100;
assign x[1143]= 32'b11110100011000101100000100010000;
assign x[1144]= 32'b11110100010010011100000100010101;
assign x[1145]= 32'b11110100001100001100000100011001;
assign x[1146]= 32'b11110100000110001100000100011110;
assign x[1147]= 32'b11110011111111111100000100100011;
assign x[1148]= 32'b11110011111001101100000100101000;
assign x[1149]= 32'b11110011110011101100000100101100;
assign x[1150]= 32'b11110011101101011100000100110001;
assign x[1151]= 32'b11110011100111001100000100110110;
assign x[1152]= 32'b11110011100001001100000100111011;
assign x[1153]= 32'b11110011011010111100000101000000;
assign x[1154]= 32'b11110011010100101100000101000101;
assign x[1155]= 32'b11110011001110101100000101001010;
assign x[1156]= 32'b11110011001000011100000101001111;
assign x[1157]= 32'b11110011000010001100000101010100;
assign x[1158]= 32'b11110010111100001100000101011001;
assign x[1159]= 32'b11110010110101111100000101011110;
assign x[1160]= 32'b11110010101111111100000101100011;
assign x[1161]= 32'b11110010101001101100000101101000;
assign x[1162]= 32'b11110010100011101100000101101110;
assign x[1163]= 32'b11110010011101011100000101110011;
assign x[1164]= 32'b11110010010111001100000101111000;
assign x[1165]= 32'b11110010010001001100000101111110;
assign x[1166]= 32'b11110010001010111100000110000011;
assign x[1167]= 32'b11110010000100111100000110001001;
assign x[1168]= 32'b11110001111110101100000110001110;
assign x[1169]= 32'b11110001111000101100000110010100;
assign x[1170]= 32'b11110001110010011100000110011001;
assign x[1171]= 32'b11110001101100011100000110011111;
assign x[1172]= 32'b11110001100110001100000110100100;
assign x[1173]= 32'b11110001100000001100000110101010;
assign x[1174]= 32'b11110001011001111100000110110000;
assign x[1175]= 32'b11110001010011111100000110110110;
assign x[1176]= 32'b11110001001101101100000110111011;
assign x[1177]= 32'b11110001000111101100000111000001;
assign x[1178]= 32'b11110001000001011100000111000111;
assign x[1179]= 32'b11110000111011011100000111001101;
assign x[1180]= 32'b11110000110101011100000111010011;
assign x[1181]= 32'b11110000101111001100000111011001;
assign x[1182]= 32'b11110000101001001100000111011111;
assign x[1183]= 32'b11110000100010111100000111100101;
assign x[1184]= 32'b11110000011100111100000111101011;
assign x[1185]= 32'b11110000010110111100000111110001;
assign x[1186]= 32'b11110000010000101100000111110111;
assign x[1187]= 32'b11110000001010101100000111111101;
assign x[1188]= 32'b11110000000100101100001000000100;
assign x[1189]= 32'b11101111111110011100001000001010;
assign x[1190]= 32'b11101111111000011100001000010000;
assign x[1191]= 32'b11101111110010011100001000010111;
assign x[1192]= 32'b11101111101100001100001000011101;
assign x[1193]= 32'b11101111100110001100001000100011;
assign x[1194]= 32'b11101111100000001100001000101010;
assign x[1195]= 32'b11101111011001111100001000110000;
assign x[1196]= 32'b11101111010011111100001000110111;
assign x[1197]= 32'b11101111001101111100001000111110;
assign x[1198]= 32'b11101111000111111100001001000100;
assign x[1199]= 32'b11101111000001101100001001001011;
assign x[1200]= 32'b11101110111011101100001001010001;
assign x[1201]= 32'b11101110110101101100001001011000;
assign x[1202]= 32'b11101110101111101100001001011111;
assign x[1203]= 32'b11101110101001101100001001100110;
assign x[1204]= 32'b11101110100011011100001001101101;
assign x[1205]= 32'b11101110011101011100001001110011;
assign x[1206]= 32'b11101110010111011100001001111010;
assign x[1207]= 32'b11101110010001011100001010000001;
assign x[1208]= 32'b11101110001011011100001010001000;
assign x[1209]= 32'b11101110000101011100001010001111;
assign x[1210]= 32'b11101101111111001100001010010110;
assign x[1211]= 32'b11101101111001001100001010011101;
assign x[1212]= 32'b11101101110011001100001010100101;
assign x[1213]= 32'b11101101101101001100001010101100;
assign x[1214]= 32'b11101101100111001100001010110011;
assign x[1215]= 32'b11101101100001001100001010111010;
assign x[1216]= 32'b11101101011011001100001011000001;
assign x[1217]= 32'b11101101010101001100001011001001;
assign x[1218]= 32'b11101101001111001100001011010000;
assign x[1219]= 32'b11101101001001001100001011011000;
assign x[1220]= 32'b11101101000011001100001011011111;
assign x[1221]= 32'b11101100111101001100001011100110;
assign x[1222]= 32'b11101100110111001100001011101110;
assign x[1223]= 32'b11101100110001001100001011110101;
assign x[1224]= 32'b11101100101011001100001011111101;
assign x[1225]= 32'b11101100100101001100001100000101;
assign x[1226]= 32'b11101100011111001100001100001100;
assign x[1227]= 32'b11101100011001001100001100010100;
assign x[1228]= 32'b11101100010011001100001100011100;
assign x[1229]= 32'b11101100001101001100001100100011;
assign x[1230]= 32'b11101100000111001100001100101011;
assign x[1231]= 32'b11101100000001011100001100110011;
assign x[1232]= 32'b11101011111011011100001100111011;
assign x[1233]= 32'b11101011110101011100001101000011;
assign x[1234]= 32'b11101011101111011100001101001011;
assign x[1235]= 32'b11101011101001011100001101010011;
assign x[1236]= 32'b11101011100011011100001101011011;
assign x[1237]= 32'b11101011011101011100001101100011;
assign x[1238]= 32'b11101011010111101100001101101011;
assign x[1239]= 32'b11101011010001101100001101110011;
assign x[1240]= 32'b11101011001011101100001101111011;
assign x[1241]= 32'b11101011000101101100001110000011;
assign x[1242]= 32'b11101010111111111100001110001100;
assign x[1243]= 32'b11101010111001111100001110010100;
assign x[1244]= 32'b11101010110011111100001110011100;
assign x[1245]= 32'b11101010101101111100001110100101;
assign x[1246]= 32'b11101010101000001100001110101101;
assign x[1247]= 32'b11101010100010001100001110110101;
assign x[1248]= 32'b11101010011100001100001110111110;
assign x[1249]= 32'b11101010010110011100001111000110;
assign x[1250]= 32'b11101010010000011100001111001111;
assign x[1251]= 32'b11101010001010011100001111010111;
assign x[1252]= 32'b11101010000100101100001111100000;
assign x[1253]= 32'b11101001111110101100001111101001;
assign x[1254]= 32'b11101001111000111100001111110001;
assign x[1255]= 32'b11101001110010111100001111111010;
assign x[1256]= 32'b11101001101101001100010000000011;
assign x[1257]= 32'b11101001100111001100010000001011;
assign x[1258]= 32'b11101001100001001100010000010100;
assign x[1259]= 32'b11101001011011011100010000011101;
assign x[1260]= 32'b11101001010101011100010000100110;
assign x[1261]= 32'b11101001001111101100010000101111;
assign x[1262]= 32'b11101001001001101100010000111000;
assign x[1263]= 32'b11101001000011111100010001000001;
assign x[1264]= 32'b11101000111101111100010001001010;
assign x[1265]= 32'b11101000111000001100010001010011;
assign x[1266]= 32'b11101000110010011100010001011100;
assign x[1267]= 32'b11101000101100011100010001100101;
assign x[1268]= 32'b11101000100110101100010001101110;
assign x[1269]= 32'b11101000100000101100010001111000;
assign x[1270]= 32'b11101000011010111100010010000001;
assign x[1271]= 32'b11101000010101001100010010001010;
assign x[1272]= 32'b11101000001111001100010010010011;
assign x[1273]= 32'b11101000001001011100010010011101;
assign x[1274]= 32'b11101000000011101100010010100110;
assign x[1275]= 32'b11100111111101101100010010110000;
assign x[1276]= 32'b11100111110111111100010010111001;
assign x[1277]= 32'b11100111110010001100010011000010;
assign x[1278]= 32'b11100111101100011100010011001100;
assign x[1279]= 32'b11100111100110011100010011010110;
assign x[1280]= 32'b11100111100000101100010011011111;
assign x[1281]= 32'b11100111011010111100010011101001;
assign x[1282]= 32'b11100111010101001100010011110010;
assign x[1283]= 32'b11100111001111011100010011111100;
assign x[1284]= 32'b11100111001001011100010100000110;
assign x[1285]= 32'b11100111000011101100010100010000;
assign x[1286]= 32'b11100110111101111100010100011010;
assign x[1287]= 32'b11100110111000001100010100100011;
assign x[1288]= 32'b11100110110010011100010100101101;
assign x[1289]= 32'b11100110101100101100010100110111;
assign x[1290]= 32'b11100110100110111100010101000001;
assign x[1291]= 32'b11100110100001001100010101001011;
assign x[1292]= 32'b11100110011011011100010101010101;
assign x[1293]= 32'b11100110010101101100010101011111;
assign x[1294]= 32'b11100110001111111100010101101001;
assign x[1295]= 32'b11100110001010001100010101110011;
assign x[1296]= 32'b11100110000100011100010101111110;
assign x[1297]= 32'b11100101111110101100010110001000;
assign x[1298]= 32'b11100101111000111100010110010010;
assign x[1299]= 32'b11100101110011001100010110011100;
assign x[1300]= 32'b11100101101101011100010110100111;
assign x[1301]= 32'b11100101100111101100010110110001;
assign x[1302]= 32'b11100101100001111100010110111011;
assign x[1303]= 32'b11100101011100001100010111000110;
assign x[1304]= 32'b11100101010110011100010111010000;
assign x[1305]= 32'b11100101010000101100010111011011;
assign x[1306]= 32'b11100101001011001100010111100101;
assign x[1307]= 32'b11100101000101011100010111110000;
assign x[1308]= 32'b11100100111111101100010111111010;
assign x[1309]= 32'b11100100111001111100011000000101;
assign x[1310]= 32'b11100100110100001100011000010000;
assign x[1311]= 32'b11100100101110101100011000011010;
assign x[1312]= 32'b11100100101000111100011000100101;
assign x[1313]= 32'b11100100100011001100011000110000;
assign x[1314]= 32'b11100100011101101100011000111011;
assign x[1315]= 32'b11100100010111111100011001000101;
assign x[1316]= 32'b11100100010010001100011001010000;
assign x[1317]= 32'b11100100001100101100011001011011;
assign x[1318]= 32'b11100100000110111100011001100110;
assign x[1319]= 32'b11100100000001001100011001110001;
assign x[1320]= 32'b11100011111011101100011001111100;
assign x[1321]= 32'b11100011110101111100011010000111;
assign x[1322]= 32'b11100011110000011100011010010010;
assign x[1323]= 32'b11100011101010101100011010011101;
assign x[1324]= 32'b11100011100101001100011010101000;
assign x[1325]= 32'b11100011011111011100011010110100;
assign x[1326]= 32'b11100011011001111100011010111111;
assign x[1327]= 32'b11100011010100001100011011001010;
assign x[1328]= 32'b11100011001110101100011011010101;
assign x[1329]= 32'b11100011001000111100011011100001;
assign x[1330]= 32'b11100011000011011100011011101100;
assign x[1331]= 32'b11100010111101101100011011110111;
assign x[1332]= 32'b11100010111000001100011100000011;
assign x[1333]= 32'b11100010110010101100011100001110;
assign x[1334]= 32'b11100010101100111100011100011010;
assign x[1335]= 32'b11100010100111011100011100100101;
assign x[1336]= 32'b11100010100001111100011100110001;
assign x[1337]= 32'b11100010011100001100011100111101;
assign x[1338]= 32'b11100010010110101100011101001000;
assign x[1339]= 32'b11100010010001001100011101010100;
assign x[1340]= 32'b11100010001011011100011101011111;
assign x[1341]= 32'b11100010000101111100011101101011;
assign x[1342]= 32'b11100010000000011100011101110111;
assign x[1343]= 32'b11100001111010111100011110000011;
assign x[1344]= 32'b11100001110101011100011110001111;
assign x[1345]= 32'b11100001101111101100011110011010;
assign x[1346]= 32'b11100001101010001100011110100110;
assign x[1347]= 32'b11100001100100101100011110110010;
assign x[1348]= 32'b11100001011111001100011110111110;
assign x[1349]= 32'b11100001011001101100011111001010;
assign x[1350]= 32'b11100001010100001100011111010110;
assign x[1351]= 32'b11100001001110101100011111100010;
assign x[1352]= 32'b11100001001001001100011111101110;
assign x[1353]= 32'b11100001000011101100011111111011;
assign x[1354]= 32'b11100000111110001100100000000111;
assign x[1355]= 32'b11100000111000101100100000010011;
assign x[1356]= 32'b11100000110011001100100000011111;
assign x[1357]= 32'b11100000101101101100100000101011;
assign x[1358]= 32'b11100000101000001100100000111000;
assign x[1359]= 32'b11100000100010101100100001000100;
assign x[1360]= 32'b11100000011101001100100001010000;
assign x[1361]= 32'b11100000010111101100100001011101;
assign x[1362]= 32'b11100000010010011100100001101001;
assign x[1363]= 32'b11100000001100111100100001110110;
assign x[1364]= 32'b11100000000111011100100010000010;
assign x[1365]= 32'b11100000000001111100100010001111;
assign x[1366]= 32'b11011111111100011100100010011011;
assign x[1367]= 32'b11011111110111001100100010101000;
assign x[1368]= 32'b11011111110001101100100010110101;
assign x[1369]= 32'b11011111101100001100100011000001;
assign x[1370]= 32'b11011111100110111100100011001110;
assign x[1371]= 32'b11011111100001011100100011011011;
assign x[1372]= 32'b11011111011011111100100011101000;
assign x[1373]= 32'b11011111010110101100100011110100;
assign x[1374]= 32'b11011111010001001100100100000001;
assign x[1375]= 32'b11011111001011111100100100001110;
assign x[1376]= 32'b11011111000110011100100100011011;
assign x[1377]= 32'b11011111000000111100100100101000;
assign x[1378]= 32'b11011110111011101100100100110101;
assign x[1379]= 32'b11011110110110001100100101000010;
assign x[1380]= 32'b11011110110000111100100101001111;
assign x[1381]= 32'b11011110101011011100100101011100;
assign x[1382]= 32'b11011110100110001100100101101001;
assign x[1383]= 32'b11011110100000111100100101110110;
assign x[1384]= 32'b11011110011011011100100110000011;
assign x[1385]= 32'b11011110010110001100100110010001;
assign x[1386]= 32'b11011110010000101100100110011110;
assign x[1387]= 32'b11011110001011011100100110101011;
assign x[1388]= 32'b11011110000110001100100110111000;
assign x[1389]= 32'b11011110000000101100100111000110;
assign x[1390]= 32'b11011101111011011100100111010011;
assign x[1391]= 32'b11011101110110001100100111100000;
assign x[1392]= 32'b11011101110000111100100111101110;
assign x[1393]= 32'b11011101101011011100100111111011;
assign x[1394]= 32'b11011101100110001100101000001001;
assign x[1395]= 32'b11011101100000111100101000010110;
assign x[1396]= 32'b11011101011011101100101000100100;
assign x[1397]= 32'b11011101010110011100101000110010;
assign x[1398]= 32'b11011101010001001100101000111111;
assign x[1399]= 32'b11011101001011101100101001001101;
assign x[1400]= 32'b11011101000110011100101001011011;
assign x[1401]= 32'b11011101000001001100101001101000;
assign x[1402]= 32'b11011100111011111100101001110110;
assign x[1403]= 32'b11011100110110101100101010000100;
assign x[1404]= 32'b11011100110001011100101010010010;
assign x[1405]= 32'b11011100101100001100101010011111;
assign x[1406]= 32'b11011100100110111100101010101101;
assign x[1407]= 32'b11011100100001101100101010111011;
assign x[1408]= 32'b11011100011100101100101011001001;
assign x[1409]= 32'b11011100010111011100101011010111;
assign x[1410]= 32'b11011100010010001100101011100101;
assign x[1411]= 32'b11011100001100111100101011110011;
assign x[1412]= 32'b11011100000111101100101100000001;
assign x[1413]= 32'b11011100000010011100101100001111;
assign x[1414]= 32'b11011011111101011100101100011110;
assign x[1415]= 32'b11011011111000001100101100101100;
assign x[1416]= 32'b11011011110010111100101100111010;
assign x[1417]= 32'b11011011101101101100101101001000;
assign x[1418]= 32'b11011011101000101100101101010110;
assign x[1419]= 32'b11011011100011011100101101100101;
assign x[1420]= 32'b11011011011110001100101101110011;
assign x[1421]= 32'b11011011011001001100101110000001;
assign x[1422]= 32'b11011011010011111100101110010000;
assign x[1423]= 32'b11011011001110111100101110011110;
assign x[1424]= 32'b11011011001001101100101110101101;
assign x[1425]= 32'b11011011000100011100101110111011;
assign x[1426]= 32'b11011010111111011100101111001010;
assign x[1427]= 32'b11011010111010001100101111011000;
assign x[1428]= 32'b11011010110101001100101111100111;
assign x[1429]= 32'b11011010101111111100101111110101;
assign x[1430]= 32'b11011010101010111100110000000100;
assign x[1431]= 32'b11011010100101111100110000010011;
assign x[1432]= 32'b11011010100000101100110000100001;
assign x[1433]= 32'b11011010011011101100110000110000;
assign x[1434]= 32'b11011010010110101100110000111111;
assign x[1435]= 32'b11011010010001011100110001001110;
assign x[1436]= 32'b11011010001100011100110001011101;
assign x[1437]= 32'b11011010000111011100110001101011;
assign x[1438]= 32'b11011010000010001100110001111010;
assign x[1439]= 32'b11011001111101001100110010001001;
assign x[1440]= 32'b11011001111000001100110010011000;
assign x[1441]= 32'b11011001110011001100110010100111;
assign x[1442]= 32'b11011001101110001100110010110110;
assign x[1443]= 32'b11011001101001001100110011000101;
assign x[1444]= 32'b11011001100011111100110011010100;
assign x[1445]= 32'b11011001011110111100110011100011;
assign x[1446]= 32'b11011001011001111100110011110011;
assign x[1447]= 32'b11011001010100111100110100000010;
assign x[1448]= 32'b11011001001111111100110100010001;
assign x[1449]= 32'b11011001001010111100110100100000;
assign x[1450]= 32'b11011001000101111100110100110000;
assign x[1451]= 32'b11011001000000111100110100111111;
assign x[1452]= 32'b11011000111011111100110101001110;
assign x[1453]= 32'b11011000110111001100110101011101;
assign x[1454]= 32'b11011000110010001100110101101101;
assign x[1455]= 32'b11011000101101001100110101111100;
assign x[1456]= 32'b11011000101000001100110110001100;
assign x[1457]= 32'b11011000100011001100110110011011;
assign x[1458]= 32'b11011000011110001100110110101011;
assign x[1459]= 32'b11011000011001011100110110111010;
assign x[1460]= 32'b11011000010100011100110111001010;
assign x[1461]= 32'b11011000001111011100110111011001;
assign x[1462]= 32'b11011000001010101100110111101001;
assign x[1463]= 32'b11011000000101101100110111111001;
assign x[1464]= 32'b11011000000000101100111000001000;
assign x[1465]= 32'b11010111111011111100111000011000;
assign x[1466]= 32'b11010111110110111100111000101000;
assign x[1467]= 32'b11010111110010001100111000111000;
assign x[1468]= 32'b11010111101101001100111001000111;
assign x[1469]= 32'b11010111101000001100111001010111;
assign x[1470]= 32'b11010111100011011100111001100111;
assign x[1471]= 32'b11010111011110101100111001110111;
assign x[1472]= 32'b11010111011001101100111010000111;
assign x[1473]= 32'b11010111010100111100111010010111;
assign x[1474]= 32'b11010111001111111100111010100111;
assign x[1475]= 32'b11010111001011001100111010110111;
assign x[1476]= 32'b11010111000110011100111011000111;
assign x[1477]= 32'b11010111000001011100111011010111;
assign x[1478]= 32'b11010110111100101100111011100111;
assign x[1479]= 32'b11010110110111111100111011110111;
assign x[1480]= 32'b11010110110010111100111100000111;
assign x[1481]= 32'b11010110101110001100111100011000;
assign x[1482]= 32'b11010110101001011100111100101000;
assign x[1483]= 32'b11010110100100101100111100111000;
assign x[1484]= 32'b11010110011111111100111101001000;
assign x[1485]= 32'b11010110011011001100111101011001;
assign x[1486]= 32'b11010110010110011100111101101001;
assign x[1487]= 32'b11010110010001011100111101111001;
assign x[1488]= 32'b11010110001100101100111110001010;
assign x[1489]= 32'b11010110000111111100111110011010;
assign x[1490]= 32'b11010110000011001100111110101011;
assign x[1491]= 32'b11010101111110011100111110111011;
assign x[1492]= 32'b11010101111001101100111111001100;
assign x[1493]= 32'b11010101110101001100111111011100;
assign x[1494]= 32'b11010101110000011100111111101101;
assign x[1495]= 32'b11010101101011101100111111111110;
assign x[1496]= 32'b11010101100110111101000000001110;
assign x[1497]= 32'b11010101100010001101000000011111;
assign x[1498]= 32'b11010101011101011101000000110000;
assign x[1499]= 32'b11010101011000111101000001000000;
assign x[1500]= 32'b11010101010100001101000001010001;
assign x[1501]= 32'b11010101001111011101000001100010;
assign x[1502]= 32'b11010101001010101101000001110011;
assign x[1503]= 32'b11010101000110001101000010000011;
assign x[1504]= 32'b11010101000001011101000010010100;
assign x[1505]= 32'b11010100111100111101000010100101;
assign x[1506]= 32'b11010100111000001101000010110110;
assign x[1507]= 32'b11010100110011011101000011000111;
assign x[1508]= 32'b11010100101110111101000011011000;
assign x[1509]= 32'b11010100101010001101000011101001;
assign x[1510]= 32'b11010100100101101101000011111010;
assign x[1511]= 32'b11010100100000111101000100001011;
assign x[1512]= 32'b11010100011100011101000100011100;
assign x[1513]= 32'b11010100010111111101000100101101;
assign x[1514]= 32'b11010100010011001101000100111110;
assign x[1515]= 32'b11010100001110101101000101010000;
assign x[1516]= 32'b11010100001010001101000101100001;
assign x[1517]= 32'b11010100000101011101000101110010;
assign x[1518]= 32'b11010100000000111101000110000011;
assign x[1519]= 32'b11010011111100011101000110010101;
assign x[1520]= 32'b11010011110111111101000110100110;
assign x[1521]= 32'b11010011110011001101000110110111;
assign x[1522]= 32'b11010011101110101101000111001001;
assign x[1523]= 32'b11010011101010001101000111011010;
assign x[1524]= 32'b11010011100101101101000111101011;
assign x[1525]= 32'b11010011100001001101000111111101;
assign x[1526]= 32'b11010011011100101101001000001110;
assign x[1527]= 32'b11010011011000001101001000100000;
assign x[1528]= 32'b11010011010011101101001000110001;
assign x[1529]= 32'b11010011001111001101001001000011;
assign x[1530]= 32'b11010011001010101101001001010101;
assign x[1531]= 32'b11010011000110001101001001100110;
assign x[1532]= 32'b11010011000001101101001001111000;
assign x[1533]= 32'b11010010111101001101001010001010;
assign x[1534]= 32'b11010010111000101101001010011011;
assign x[1535]= 32'b11010010110100011101001010101101;
assign x[1536]= 32'b11010010101111111101001010111111;
assign x[1537]= 32'b11010010101011011101001011010001;
assign x[1538]= 32'b11010010100110111101001011100010;
assign x[1539]= 32'b11010010100010101101001011110100;
assign x[1540]= 32'b11010010011110001101001100000110;
assign x[1541]= 32'b11010010011001101101001100011000;
assign x[1542]= 32'b11010010010101011101001100101010;
assign x[1543]= 32'b11010010010000111101001100111100;
assign x[1544]= 32'b11010010001100011101001101001110;
assign x[1545]= 32'b11010010001000001101001101100000;
assign x[1546]= 32'b11010010000011101101001101110010;
assign x[1547]= 32'b11010001111111011101001110000100;
assign x[1548]= 32'b11010001111010111101001110010110;
assign x[1549]= 32'b11010001110110101101001110101000;
assign x[1550]= 32'b11010001110010011101001110111010;
assign x[1551]= 32'b11010001101101111101001111001100;
assign x[1552]= 32'b11010001101001101101001111011111;
assign x[1553]= 32'b11010001100101011101001111110001;
assign x[1554]= 32'b11010001100000111101010000000011;
assign x[1555]= 32'b11010001011100101101010000010101;
assign x[1556]= 32'b11010001011000011101010000101000;
assign x[1557]= 32'b11010001010100001101010000111010;
assign x[1558]= 32'b11010001001111101101010001001100;
assign x[1559]= 32'b11010001001011011101010001011111;
assign x[1560]= 32'b11010001000111001101010001110001;
assign x[1561]= 32'b11010001000010111101010010000011;
assign x[1562]= 32'b11010000111110101101010010010110;
assign x[1563]= 32'b11010000111010011101010010101000;
assign x[1564]= 32'b11010000110110001101010010111011;
assign x[1565]= 32'b11010000110001111101010011001101;
assign x[1566]= 32'b11010000101101101101010011100000;
assign x[1567]= 32'b11010000101001011101010011110011;
assign x[1568]= 32'b11010000100101001101010100000101;
assign x[1569]= 32'b11010000100000111101010100011000;
assign x[1570]= 32'b11010000011100111101010100101010;
assign x[1571]= 32'b11010000011000101101010100111101;
assign x[1572]= 32'b11010000010100011101010101010000;
assign x[1573]= 32'b11010000010000001101010101100011;
assign x[1574]= 32'b11010000001100001101010101110101;
assign x[1575]= 32'b11010000000111111101010110001000;
assign x[1576]= 32'b11010000000011101101010110011011;
assign x[1577]= 32'b11001111111111101101010110101110;
assign x[1578]= 32'b11001111111011011101010111000001;
assign x[1579]= 32'b11001111110111001101010111010100;
assign x[1580]= 32'b11001111110011001101010111100110;
assign x[1581]= 32'b11001111101110111101010111111001;
assign x[1582]= 32'b11001111101010111101011000001100;
assign x[1583]= 32'b11001111100110101101011000011111;
assign x[1584]= 32'b11001111100010101101011000110010;
assign x[1585]= 32'b11001111011110011101011001000101;
assign x[1586]= 32'b11001111011010011101011001011001;
assign x[1587]= 32'b11001111010110011101011001101100;
assign x[1588]= 32'b11001111010010001101011001111111;
assign x[1589]= 32'b11001111001110001101011010010010;
assign x[1590]= 32'b11001111001010001101011010100101;
assign x[1591]= 32'b11001111000110001101011010111000;
assign x[1592]= 32'b11001111000001111101011011001011;
assign x[1593]= 32'b11001110111101111101011011011111;
assign x[1594]= 32'b11001110111001111101011011110010;
assign x[1595]= 32'b11001110110101111101011100000101;
assign x[1596]= 32'b11001110110001111101011100011001;
assign x[1597]= 32'b11001110101101111101011100101100;
assign x[1598]= 32'b11001110101001111101011100111111;
assign x[1599]= 32'b11001110100101111101011101010011;
assign x[1600]= 32'b11001110100001111101011101100110;
assign x[1601]= 32'b11001110011101111101011101111010;
assign x[1602]= 32'b11001110011001111101011110001101;
assign x[1603]= 32'b11001110010101111101011110100000;
assign x[1604]= 32'b11001110010001111101011110110100;
assign x[1605]= 32'b11001110001110001101011111001000;
assign x[1606]= 32'b11001110001010001101011111011011;
assign x[1607]= 32'b11001110000110001101011111101111;
assign x[1608]= 32'b11001110000010001101100000000010;
assign x[1609]= 32'b11001101111110011101100000010110;
assign x[1610]= 32'b11001101111010011101100000101010;
assign x[1611]= 32'b11001101110110011101100000111101;
assign x[1612]= 32'b11001101110010101101100001010001;
assign x[1613]= 32'b11001101101110101101100001100101;
assign x[1614]= 32'b11001101101010111101100001111000;
assign x[1615]= 32'b11001101100110111101100010001100;
assign x[1616]= 32'b11001101100011001101100010100000;
assign x[1617]= 32'b11001101011111001101100010110100;
assign x[1618]= 32'b11001101011011011101100011001000;
assign x[1619]= 32'b11001101010111011101100011011100;
assign x[1620]= 32'b11001101010011101101100011101111;
assign x[1621]= 32'b11001101001111111101100100000011;
assign x[1622]= 32'b11001101001100001101100100010111;
assign x[1623]= 32'b11001101001000001101100100101011;
assign x[1624]= 32'b11001101000100011101100100111111;
assign x[1625]= 32'b11001101000000101101100101010011;
assign x[1626]= 32'b11001100111100111101100101100111;
assign x[1627]= 32'b11001100111000111101100101111011;
assign x[1628]= 32'b11001100110101001101100110001111;
assign x[1629]= 32'b11001100110001011101100110100100;
assign x[1630]= 32'b11001100101101101101100110111000;
assign x[1631]= 32'b11001100101001111101100111001100;
assign x[1632]= 32'b11001100100110001101100111100000;
assign x[1633]= 32'b11001100100010011101100111110100;
assign x[1634]= 32'b11001100011110101101101000001000;
assign x[1635]= 32'b11001100011010111101101000011101;
assign x[1636]= 32'b11001100010111011101101000110001;
assign x[1637]= 32'b11001100010011101101101001000101;
assign x[1638]= 32'b11001100001111111101101001011010;
assign x[1639]= 32'b11001100001100001101101001101110;
assign x[1640]= 32'b11001100001000011101101010000010;
assign x[1641]= 32'b11001100000100111101101010010111;
assign x[1642]= 32'b11001100000001001101101010101011;
assign x[1643]= 32'b11001011111101011101101010111111;
assign x[1644]= 32'b11001011111001111101101011010100;
assign x[1645]= 32'b11001011110110001101101011101000;
assign x[1646]= 32'b11001011110010101101101011111101;
assign x[1647]= 32'b11001011101110111101101100010001;
assign x[1648]= 32'b11001011101011011101101100100110;
assign x[1649]= 32'b11001011100111101101101100111011;
assign x[1650]= 32'b11001011100100001101101101001111;
assign x[1651]= 32'b11001011100000011101101101100100;
assign x[1652]= 32'b11001011011100111101101101111000;
assign x[1653]= 32'b11001011011001011101101110001101;
assign x[1654]= 32'b11001011010101101101101110100010;
assign x[1655]= 32'b11001011010010001101101110110110;
assign x[1656]= 32'b11001011001110101101101111001011;
assign x[1657]= 32'b11001011001011001101101111100000;
assign x[1658]= 32'b11001011000111101101101111110101;
assign x[1659]= 32'b11001011000011111101110000001001;
assign x[1660]= 32'b11001011000000011101110000011110;
assign x[1661]= 32'b11001010111100111101110000110011;
assign x[1662]= 32'b11001010111001011101110001001000;
assign x[1663]= 32'b11001010110101111101110001011101;
assign x[1664]= 32'b11001010110010011101110001110010;
assign x[1665]= 32'b11001010101110111101110010000110;
assign x[1666]= 32'b11001010101011011101110010011011;
assign x[1667]= 32'b11001010100111111101110010110000;
assign x[1668]= 32'b11001010100100101101110011000101;
assign x[1669]= 32'b11001010100001001101110011011010;
assign x[1670]= 32'b11001010011101101101110011101111;
assign x[1671]= 32'b11001010011010001101110100000100;
assign x[1672]= 32'b11001010010110111101110100011001;
assign x[1673]= 32'b11001010010011011101110100101110;
assign x[1674]= 32'b11001010001111111101110101000100;
assign x[1675]= 32'b11001010001100101101110101011001;
assign x[1676]= 32'b11001010001001001101110101101110;
assign x[1677]= 32'b11001010000101101101110110000011;
assign x[1678]= 32'b11001010000010011101110110011000;
assign x[1679]= 32'b11001001111110111101110110101101;
assign x[1680]= 32'b11001001111011101101110111000011;
assign x[1681]= 32'b11001001111000001101110111011000;
assign x[1682]= 32'b11001001110100111101110111101101;
assign x[1683]= 32'b11001001110001101101111000000010;
assign x[1684]= 32'b11001001101110001101111000011000;
assign x[1685]= 32'b11001001101010111101111000101101;
assign x[1686]= 32'b11001001100111101101111001000010;
assign x[1687]= 32'b11001001100100011101111001011000;
assign x[1688]= 32'b11001001100000111101111001101101;
assign x[1689]= 32'b11001001011101101101111010000011;
assign x[1690]= 32'b11001001011010011101111010011000;
assign x[1691]= 32'b11001001010111001101111010101101;
assign x[1692]= 32'b11001001010011111101111011000011;
assign x[1693]= 32'b11001001010000101101111011011000;
assign x[1694]= 32'b11001001001101011101111011101110;
assign x[1695]= 32'b11001001001010001101111100000011;
assign x[1696]= 32'b11001001000110111101111100011001;
assign x[1697]= 32'b11001001000011101101111100101111;
assign x[1698]= 32'b11001001000000011101111101000100;
assign x[1699]= 32'b11001000111101001101111101011010;
assign x[1700]= 32'b11001000111010001101111101101111;
assign x[1701]= 32'b11001000110110111101111110000101;
assign x[1702]= 32'b11001000110011101101111110011011;
assign x[1703]= 32'b11001000110000011101111110110000;
assign x[1704]= 32'b11001000101101011101111111000110;
assign x[1705]= 32'b11001000101010001101111111011100;
assign x[1706]= 32'b11001000100110111101111111110001;
assign x[1707]= 32'b11001000100011111110000000000111;
assign x[1708]= 32'b11001000100000101110000000011101;
assign x[1709]= 32'b11001000011101101110000000110011;
assign x[1710]= 32'b11001000011010011110000001001001;
assign x[1711]= 32'b11001000010111011110000001011110;
assign x[1712]= 32'b11001000010100001110000001110100;
assign x[1713]= 32'b11001000010001001110000010001010;
assign x[1714]= 32'b11001000001110001110000010100000;
assign x[1715]= 32'b11001000001010111110000010110110;
assign x[1716]= 32'b11001000000111111110000011001100;
assign x[1717]= 32'b11001000000100111110000011100010;
assign x[1718]= 32'b11001000000001111110000011111000;
assign x[1719]= 32'b11000111111110111110000100001110;
assign x[1720]= 32'b11000111111011101110000100100100;
assign x[1721]= 32'b11000111111000101110000100111010;
assign x[1722]= 32'b11000111110101101110000101010000;
assign x[1723]= 32'b11000111110010101110000101100110;
assign x[1724]= 32'b11000111101111101110000101111100;
assign x[1725]= 32'b11000111101100101110000110010010;
assign x[1726]= 32'b11000111101001101110000110101000;
assign x[1727]= 32'b11000111100110101110000110111110;
assign x[1728]= 32'b11000111100011111110000111010101;
assign x[1729]= 32'b11000111100000111110000111101011;
assign x[1730]= 32'b11000111011101111110001000000001;
assign x[1731]= 32'b11000111011010111110001000010111;
assign x[1732]= 32'b11000111010111111110001000101101;
assign x[1733]= 32'b11000111010101001110001001000100;
assign x[1734]= 32'b11000111010010001110001001011010;
assign x[1735]= 32'b11000111001111011110001001110000;
assign x[1736]= 32'b11000111001100011110001010000111;
assign x[1737]= 32'b11000111001001011110001010011101;
assign x[1738]= 32'b11000111000110101110001010110011;
assign x[1739]= 32'b11000111000011101110001011001010;
assign x[1740]= 32'b11000111000000111110001011100000;
assign x[1741]= 32'b11000110111101111110001011110110;
assign x[1742]= 32'b11000110111011001110001100001101;
assign x[1743]= 32'b11000110111000011110001100100011;
assign x[1744]= 32'b11000110110101011110001100111010;
assign x[1745]= 32'b11000110110010101110001101010000;
assign x[1746]= 32'b11000110101111111110001101100111;
assign x[1747]= 32'b11000110101101001110001101111101;
assign x[1748]= 32'b11000110101010001110001110010100;
assign x[1749]= 32'b11000110100111011110001110101010;
assign x[1750]= 32'b11000110100100101110001111000001;
assign x[1751]= 32'b11000110100001111110001111010111;
assign x[1752]= 32'b11000110011111001110001111101110;
assign x[1753]= 32'b11000110011100011110010000000100;
assign x[1754]= 32'b11000110011001101110010000011011;
assign x[1755]= 32'b11000110010110111110010000110010;
assign x[1756]= 32'b11000110010100001110010001001000;
assign x[1757]= 32'b11000110010001011110010001011111;
assign x[1758]= 32'b11000110001110111110010001110110;
assign x[1759]= 32'b11000110001100001110010010001100;
assign x[1760]= 32'b11000110001001011110010010100011;
assign x[1761]= 32'b11000110000110101110010010111010;
assign x[1762]= 32'b11000110000100001110010011010000;
assign x[1763]= 32'b11000110000001011110010011100111;
assign x[1764]= 32'b11000101111110101110010011111110;
assign x[1765]= 32'b11000101111100001110010100010101;
assign x[1766]= 32'b11000101111001011110010100101100;
assign x[1767]= 32'b11000101110110111110010101000010;
assign x[1768]= 32'b11000101110100001110010101011001;
assign x[1769]= 32'b11000101110001101110010101110000;
assign x[1770]= 32'b11000101101110111110010110000111;
assign x[1771]= 32'b11000101101100011110010110011110;
assign x[1772]= 32'b11000101101001111110010110110101;
assign x[1773]= 32'b11000101100111001110010111001100;
assign x[1774]= 32'b11000101100100101110010111100011;
assign x[1775]= 32'b11000101100010001110010111111010;
assign x[1776]= 32'b11000101011111101110011000010001;
assign x[1777]= 32'b11000101011100111110011000101000;
assign x[1778]= 32'b11000101011010011110011000111111;
assign x[1779]= 32'b11000101010111111110011001010110;
assign x[1780]= 32'b11000101010101011110011001101101;
assign x[1781]= 32'b11000101010010111110011010000100;
assign x[1782]= 32'b11000101010000011110011010011011;
assign x[1783]= 32'b11000101001101111110011010110010;
assign x[1784]= 32'b11000101001011011110011011001001;
assign x[1785]= 32'b11000101001000111110011011100000;
assign x[1786]= 32'b11000101000110101110011011110111;
assign x[1787]= 32'b11000101000100001110011100001110;
assign x[1788]= 32'b11000101000001101110011100100101;
assign x[1789]= 32'b11000100111111001110011100111101;
assign x[1790]= 32'b11000100111100101110011101010100;
assign x[1791]= 32'b11000100111010011110011101101011;
assign x[1792]= 32'b11000100110111111110011110000010;
assign x[1793]= 32'b11000100110101101110011110011001;
assign x[1794]= 32'b11000100110011001110011110110001;
assign x[1795]= 32'b11000100110000101110011111001000;
assign x[1796]= 32'b11000100101110011110011111011111;
assign x[1797]= 32'b11000100101100001110011111110110;
assign x[1798]= 32'b11000100101001101110100000001110;
assign x[1799]= 32'b11000100100111011110100000100101;
assign x[1800]= 32'b11000100100100111110100000111100;
assign x[1801]= 32'b11000100100010101110100001010100;
assign x[1802]= 32'b11000100100000011110100001101011;
assign x[1803]= 32'b11000100011110001110100010000010;
assign x[1804]= 32'b11000100011011101110100010011010;
assign x[1805]= 32'b11000100011001011110100010110001;
assign x[1806]= 32'b11000100010111001110100011001001;
assign x[1807]= 32'b11000100010100111110100011100000;
assign x[1808]= 32'b11000100010010101110100011110111;
assign x[1809]= 32'b11000100010000011110100100001111;
assign x[1810]= 32'b11000100001110001110100100100110;
assign x[1811]= 32'b11000100001011111110100100111110;
assign x[1812]= 32'b11000100001001101110100101010101;
assign x[1813]= 32'b11000100000111011110100101101101;
assign x[1814]= 32'b11000100000101001110100110000100;
assign x[1815]= 32'b11000100000010111110100110011100;
assign x[1816]= 32'b11000100000000111110100110110100;
assign x[1817]= 32'b11000011111110101110100111001011;
assign x[1818]= 32'b11000011111100011110100111100011;
assign x[1819]= 32'b11000011111010011110100111111010;
assign x[1820]= 32'b11000011111000001110101000010010;
assign x[1821]= 32'b11000011110101111110101000101001;
assign x[1822]= 32'b11000011110011111110101001000001;
assign x[1823]= 32'b11000011110001101110101001011001;
assign x[1824]= 32'b11000011101111101110101001110000;
assign x[1825]= 32'b11000011101101011110101010001000;
assign x[1826]= 32'b11000011101011011110101010100000;
assign x[1827]= 32'b11000011101001011110101010110111;
assign x[1828]= 32'b11000011100111001110101011001111;
assign x[1829]= 32'b11000011100101001110101011100111;
assign x[1830]= 32'b11000011100011001110101011111111;
assign x[1831]= 32'b11000011100000111110101100010110;
assign x[1832]= 32'b11000011011110111110101100101110;
assign x[1833]= 32'b11000011011100111110101101000110;
assign x[1834]= 32'b11000011011010111110101101011110;
assign x[1835]= 32'b11000011011000111110101101110101;
assign x[1836]= 32'b11000011010110111110101110001101;
assign x[1837]= 32'b11000011010100111110101110100101;
assign x[1838]= 32'b11000011010010111110101110111101;
assign x[1839]= 32'b11000011010000111110101111010101;
assign x[1840]= 32'b11000011001110111110101111101101;
assign x[1841]= 32'b11000011001100111110110000000101;
assign x[1842]= 32'b11000011001010111110110000011100;
assign x[1843]= 32'b11000011001000111110110000110100;
assign x[1844]= 32'b11000011000111001110110001001100;
assign x[1845]= 32'b11000011000101001110110001100100;
assign x[1846]= 32'b11000011000011001110110001111100;
assign x[1847]= 32'b11000011000001011110110010010100;
assign x[1848]= 32'b11000010111111011110110010101100;
assign x[1849]= 32'b11000010111101011110110011000100;
assign x[1850]= 32'b11000010111011101110110011011100;
assign x[1851]= 32'b11000010111001101110110011110100;
assign x[1852]= 32'b11000010110111111110110100001100;
assign x[1853]= 32'b11000010110110001110110100100100;
assign x[1854]= 32'b11000010110100001110110100111100;
assign x[1855]= 32'b11000010110010011110110101010100;
assign x[1856]= 32'b11000010110000011110110101101100;
assign x[1857]= 32'b11000010101110101110110110000100;
assign x[1858]= 32'b11000010101100111110110110011100;
assign x[1859]= 32'b11000010101011001110110110110100;
assign x[1860]= 32'b11000010101001011110110111001100;
assign x[1861]= 32'b11000010100111011110110111100100;
assign x[1862]= 32'b11000010100101101110110111111100;
assign x[1863]= 32'b11000010100011111110111000010101;
assign x[1864]= 32'b11000010100010001110111000101101;
assign x[1865]= 32'b11000010100000011110111001000101;
assign x[1866]= 32'b11000010011110101110111001011101;
assign x[1867]= 32'b11000010011100111110111001110101;
assign x[1868]= 32'b11000010011011011110111010001101;
assign x[1869]= 32'b11000010011001101110111010100110;
assign x[1870]= 32'b11000010010111111110111010111110;
assign x[1871]= 32'b11000010010110001110111011010110;
assign x[1872]= 32'b11000010010100011110111011101110;
assign x[1873]= 32'b11000010010010111110111100000110;
assign x[1874]= 32'b11000010010001001110111100011111;
assign x[1875]= 32'b11000010001111101110111100110111;
assign x[1876]= 32'b11000010001101111110111101001111;
assign x[1877]= 32'b11000010001100001110111101100111;
assign x[1878]= 32'b11000010001010101110111110000000;
assign x[1879]= 32'b11000010001000111110111110011000;
assign x[1880]= 32'b11000010000111011110111110110000;
assign x[1881]= 32'b11000010000101111110111111001001;
assign x[1882]= 32'b11000010000100001110111111100001;
assign x[1883]= 32'b11000010000010101110111111111001;
assign x[1884]= 32'b11000010000001001111000000010010;
assign x[1885]= 32'b11000001111111011111000000101010;
assign x[1886]= 32'b11000001111101111111000001000010;
assign x[1887]= 32'b11000001111100011111000001011011;
assign x[1888]= 32'b11000001111010111111000001110011;
assign x[1889]= 32'b11000001111001011111000010001011;
assign x[1890]= 32'b11000001110111111111000010100100;
assign x[1891]= 32'b11000001110110011111000010111100;
assign x[1892]= 32'b11000001110100111111000011010101;
assign x[1893]= 32'b11000001110011011111000011101101;
assign x[1894]= 32'b11000001110001111111000100000101;
assign x[1895]= 32'b11000001110000011111000100011110;
assign x[1896]= 32'b11000001101110111111000100110110;
assign x[1897]= 32'b11000001101101101111000101001111;
assign x[1898]= 32'b11000001101100001111000101100111;
assign x[1899]= 32'b11000001101010101111000110000000;
assign x[1900]= 32'b11000001101001001111000110011000;
assign x[1901]= 32'b11000001100111111111000110110001;
assign x[1902]= 32'b11000001100110011111000111001001;
assign x[1903]= 32'b11000001100101001111000111100010;
assign x[1904]= 32'b11000001100011101111000111111010;
assign x[1905]= 32'b11000001100010011111001000010011;
assign x[1906]= 32'b11000001100000111111001000101011;
assign x[1907]= 32'b11000001011111101111001001000100;
assign x[1908]= 32'b11000001011110001111001001011100;
assign x[1909]= 32'b11000001011100111111001001110101;
assign x[1910]= 32'b11000001011011101111001010001110;
assign x[1911]= 32'b11000001011010001111001010100110;
assign x[1912]= 32'b11000001011000111111001010111111;
assign x[1913]= 32'b11000001010111101111001011010111;
assign x[1914]= 32'b11000001010110011111001011110000;
assign x[1915]= 32'b11000001010101001111001100001000;
assign x[1916]= 32'b11000001010011111111001100100001;
assign x[1917]= 32'b11000001010010101111001100111010;
assign x[1918]= 32'b11000001010001011111001101010010;
assign x[1919]= 32'b11000001010000001111001101101011;
assign x[1920]= 32'b11000001001110111111001110000100;
assign x[1921]= 32'b11000001001101101111001110011100;
assign x[1922]= 32'b11000001001100011111001110110101;
assign x[1923]= 32'b11000001001011001111001111001110;
assign x[1924]= 32'b11000001001010001111001111100110;
assign x[1925]= 32'b11000001001000111111001111111111;
assign x[1926]= 32'b11000001000111101111010000011000;
assign x[1927]= 32'b11000001000110011111010000110000;
assign x[1928]= 32'b11000001000101011111010001001001;
assign x[1929]= 32'b11000001000100001111010001100010;
assign x[1930]= 32'b11000001000011001111010001111011;
assign x[1931]= 32'b11000001000001111111010010010011;
assign x[1932]= 32'b11000001000000111111010010101100;
assign x[1933]= 32'b11000000111111101111010011000101;
assign x[1934]= 32'b11000000111110101111010011011101;
assign x[1935]= 32'b11000000111101101111010011110110;
assign x[1936]= 32'b11000000111100011111010100001111;
assign x[1937]= 32'b11000000111011011111010100101000;
assign x[1938]= 32'b11000000111010011111010101000000;
assign x[1939]= 32'b11000000111001001111010101011001;
assign x[1940]= 32'b11000000111000001111010101110010;
assign x[1941]= 32'b11000000110111001111010110001011;
assign x[1942]= 32'b11000000110110001111010110100100;
assign x[1943]= 32'b11000000110101001111010110111100;
assign x[1944]= 32'b11000000110100001111010111010101;
assign x[1945]= 32'b11000000110011001111010111101110;
assign x[1946]= 32'b11000000110010001111011000000111;
assign x[1947]= 32'b11000000110001001111011000100000;
assign x[1948]= 32'b11000000110000001111011000111001;
assign x[1949]= 32'b11000000101111011111011001010001;
assign x[1950]= 32'b11000000101110011111011001101010;
assign x[1951]= 32'b11000000101101011111011010000011;
assign x[1952]= 32'b11000000101100011111011010011100;
assign x[1953]= 32'b11000000101011101111011010110101;
assign x[1954]= 32'b11000000101010101111011011001110;
assign x[1955]= 32'b11000000101001101111011011100111;
assign x[1956]= 32'b11000000101000111111011011111111;
assign x[1957]= 32'b11000000100111111111011100011000;
assign x[1958]= 32'b11000000100111001111011100110001;
assign x[1959]= 32'b11000000100110001111011101001010;
assign x[1960]= 32'b11000000100101011111011101100011;
assign x[1961]= 32'b11000000100100101111011101111100;
assign x[1962]= 32'b11000000100011101111011110010101;
assign x[1963]= 32'b11000000100010111111011110101110;
assign x[1964]= 32'b11000000100010001111011111000111;
assign x[1965]= 32'b11000000100001011111011111100000;
assign x[1966]= 32'b11000000100000011111011111111001;
assign x[1967]= 32'b11000000011111101111100000010001;
assign x[1968]= 32'b11000000011110111111100000101010;
assign x[1969]= 32'b11000000011110001111100001000011;
assign x[1970]= 32'b11000000011101011111100001011100;
assign x[1971]= 32'b11000000011100101111100001110101;
assign x[1972]= 32'b11000000011011111111100010001110;
assign x[1973]= 32'b11000000011011001111100010100111;
assign x[1974]= 32'b11000000011010011111100011000000;
assign x[1975]= 32'b11000000011001111111100011011001;
assign x[1976]= 32'b11000000011001001111100011110010;
assign x[1977]= 32'b11000000011000011111100100001011;
assign x[1978]= 32'b11000000010111101111100100100100;
assign x[1979]= 32'b11000000010111001111100100111101;
assign x[1980]= 32'b11000000010110011111100101010110;
assign x[1981]= 32'b11000000010101101111100101101111;
assign x[1982]= 32'b11000000010101001111100110001000;
assign x[1983]= 32'b11000000010100011111100110100001;
assign x[1984]= 32'b11000000010011111111100110111010;
assign x[1985]= 32'b11000000010011001111100111010011;
assign x[1986]= 32'b11000000010010101111100111101100;
assign x[1987]= 32'b11000000010010001111101000000101;
assign x[1988]= 32'b11000000010001011111101000011110;
assign x[1989]= 32'b11000000010000111111101000110111;
assign x[1990]= 32'b11000000010000011111101001010000;
assign x[1991]= 32'b11000000001111111111101001101001;
assign x[1992]= 32'b11000000001111001111101010000010;
assign x[1993]= 32'b11000000001110101111101010011011;
assign x[1994]= 32'b11000000001110001111101010110100;
assign x[1995]= 32'b11000000001101101111101011001101;
assign x[1996]= 32'b11000000001101001111101011100110;
assign x[1997]= 32'b11000000001100101111101100000000;
assign x[1998]= 32'b11000000001100001111101100011001;
assign x[1999]= 32'b11000000001011101111101100110010;
assign x[2000]= 32'b11000000001011001111101101001011;
assign x[2001]= 32'b11000000001010111111101101100100;
assign x[2002]= 32'b11000000001010011111101101111101;
assign x[2003]= 32'b11000000001001111111101110010110;
assign x[2004]= 32'b11000000001001011111101110101111;
assign x[2005]= 32'b11000000001001001111101111001000;
assign x[2006]= 32'b11000000001000101111101111100001;
assign x[2007]= 32'b11000000001000001111101111111010;
assign x[2008]= 32'b11000000000111111111110000010011;
assign x[2009]= 32'b11000000000111011111110000101100;
assign x[2010]= 32'b11000000000111001111110001000101;
assign x[2011]= 32'b11000000000110101111110001011111;
assign x[2012]= 32'b11000000000110011111110001111000;
assign x[2013]= 32'b11000000000110001111110010010001;
assign x[2014]= 32'b11000000000101101111110010101010;
assign x[2015]= 32'b11000000000101011111110011000011;
assign x[2016]= 32'b11000000000101001111110011011100;
assign x[2017]= 32'b11000000000100111111110011110101;
assign x[2018]= 32'b11000000000100011111110100001110;
assign x[2019]= 32'b11000000000100001111110100100111;
assign x[2020]= 32'b11000000000011111111110101000000;
assign x[2021]= 32'b11000000000011101111110101011010;
assign x[2022]= 32'b11000000000011011111110101110011;
assign x[2023]= 32'b11000000000011001111110110001100;
assign x[2024]= 32'b11000000000010111111110110100101;
assign x[2025]= 32'b11000000000010101111110110111110;
assign x[2026]= 32'b11000000000010011111110111010111;
assign x[2027]= 32'b11000000000010011111110111110000;
assign x[2028]= 32'b11000000000010001111111000001001;
assign x[2029]= 32'b11000000000001111111111000100011;
assign x[2030]= 32'b11000000000001101111111000111100;
assign x[2031]= 32'b11000000000001101111111001010101;
assign x[2032]= 32'b11000000000001011111111001101110;
assign x[2033]= 32'b11000000000001001111111010000111;
assign x[2034]= 32'b11000000000001001111111010100000;
assign x[2035]= 32'b11000000000000111111111010111001;
assign x[2036]= 32'b11000000000000111111111011010010;
assign x[2037]= 32'b11000000000000101111111011101100;
assign x[2038]= 32'b11000000000000101111111100000101;
assign x[2039]= 32'b11000000000000101111111100011110;
assign x[2040]= 32'b11000000000000011111111100110111;
assign x[2041]= 32'b11000000000000011111111101010000;
assign x[2042]= 32'b11000000000000011111111101101001;
assign x[2043]= 32'b11000000000000001111111110000010;
assign x[2044]= 32'b11000000000000001111111110011011;
assign x[2045]= 32'b11000000000000001111111110110101;
assign x[2046]= 32'b11000000000000001111111111001110;
assign x[2047]= 32'b11000000000000001111111111100111;
assign x[2048]= 32'b11000000000000001111111111111111;
assign x[2049]= 32'b11000000000000000000000000011001;
assign x[2050]= 32'b11000000000000000000000000110010;
assign x[2051]= 32'b11000000000000000000000001001011;
assign x[2052]= 32'b11000000000000000000000001100100;
assign x[2053]= 32'b11000000000000000000000001111101;
assign x[2054]= 32'b11000000000000010000000010010110;
assign x[2055]= 32'b11000000000000010000000010101111;
assign x[2056]= 32'b11000000000000010000000011001001;
assign x[2057]= 32'b11000000000000100000000011100010;
assign x[2058]= 32'b11000000000000100000000011111011;
assign x[2059]= 32'b11000000000000100000000100010100;
assign x[2060]= 32'b11000000000000110000000100101101;
assign x[2061]= 32'b11000000000000110000000101000110;
assign x[2062]= 32'b11000000000001000000000101011111;
assign x[2063]= 32'b11000000000001000000000101111000;
assign x[2064]= 32'b11000000000001010000000110010010;
assign x[2065]= 32'b11000000000001100000000110101011;
assign x[2066]= 32'b11000000000001100000000111000100;
assign x[2067]= 32'b11000000000001110000000111011101;
assign x[2068]= 32'b11000000000010000000000111110110;
assign x[2069]= 32'b11000000000010010000001000001111;
assign x[2070]= 32'b11000000000010010000001000101000;
assign x[2071]= 32'b11000000000010100000001001000001;
assign x[2072]= 32'b11000000000010110000001001011011;
assign x[2073]= 32'b11000000000011000000001001110100;
assign x[2074]= 32'b11000000000011010000001010001101;
assign x[2075]= 32'b11000000000011100000001010100110;
assign x[2076]= 32'b11000000000011110000001010111111;
assign x[2077]= 32'b11000000000100000000001011011000;
assign x[2078]= 32'b11000000000100010000001011110001;
assign x[2079]= 32'b11000000000100110000001100001010;
assign x[2080]= 32'b11000000000101000000001100100011;
assign x[2081]= 32'b11000000000101010000001100111101;
assign x[2082]= 32'b11000000000101100000001101010110;
assign x[2083]= 32'b11000000000110000000001101101111;
assign x[2084]= 32'b11000000000110010000001110001000;
assign x[2085]= 32'b11000000000110100000001110100001;
assign x[2086]= 32'b11000000000111000000001110111010;
assign x[2087]= 32'b11000000000111010000001111010011;
assign x[2088]= 32'b11000000000111110000001111101100;
assign x[2089]= 32'b11000000001000000000010000000101;
assign x[2090]= 32'b11000000001000100000010000011110;
assign x[2091]= 32'b11000000001001000000010000110111;
assign x[2092]= 32'b11000000001001010000010001010001;
assign x[2093]= 32'b11000000001001110000010001101010;
assign x[2094]= 32'b11000000001010010000010010000011;
assign x[2095]= 32'b11000000001010110000010010011100;
assign x[2096]= 32'b11000000001011000000010010110101;
assign x[2097]= 32'b11000000001011100000010011001110;
assign x[2098]= 32'b11000000001100000000010011100111;
assign x[2099]= 32'b11000000001100100000010100000000;
assign x[2100]= 32'b11000000001101000000010100011001;
assign x[2101]= 32'b11000000001101100000010100110010;
assign x[2102]= 32'b11000000001110000000010101001011;
assign x[2103]= 32'b11000000001110100000010101100100;
assign x[2104]= 32'b11000000001111000000010101111101;
assign x[2105]= 32'b11000000001111110000010110010110;
assign x[2106]= 32'b11000000010000010000010110101111;
assign x[2107]= 32'b11000000010000110000010111001000;
assign x[2108]= 32'b11000000010001010000010111100001;
assign x[2109]= 32'b11000000010010000000010111111010;
assign x[2110]= 32'b11000000010010100000011000010011;
assign x[2111]= 32'b11000000010011000000011000101100;
assign x[2112]= 32'b11000000010011110000011001000101;
assign x[2113]= 32'b11000000010100010000011001011110;
assign x[2114]= 32'b11000000010101000000011001110111;
assign x[2115]= 32'b11000000010101100000011010010000;
assign x[2116]= 32'b11000000010110010000011010101001;
assign x[2117]= 32'b11000000010111000000011011000010;
assign x[2118]= 32'b11000000010111100000011011011011;
assign x[2119]= 32'b11000000011000010000011011110100;
assign x[2120]= 32'b11000000011001000000011100001101;
assign x[2121]= 32'b11000000011001110000011100100110;
assign x[2122]= 32'b11000000011010010000011100111111;
assign x[2123]= 32'b11000000011011000000011101011000;
assign x[2124]= 32'b11000000011011110000011101110001;
assign x[2125]= 32'b11000000011100100000011110001010;
assign x[2126]= 32'b11000000011101010000011110100011;
assign x[2127]= 32'b11000000011110000000011110111100;
assign x[2128]= 32'b11000000011110110000011111010101;
assign x[2129]= 32'b11000000011111100000011111101110;
assign x[2130]= 32'b11000000100000010000100000000111;
assign x[2131]= 32'b11000000100001010000100000100000;
assign x[2132]= 32'b11000000100010000000100000111001;
assign x[2133]= 32'b11000000100010110000100001010010;
assign x[2134]= 32'b11000000100011100000100001101011;
assign x[2135]= 32'b11000000100100100000100010000100;
assign x[2136]= 32'b11000000100101010000100010011100;
assign x[2137]= 32'b11000000100110000000100010110101;
assign x[2138]= 32'b11000000100111000000100011001110;
assign x[2139]= 32'b11000000100111110000100011100111;
assign x[2140]= 32'b11000000101000110000100100000000;
assign x[2141]= 32'b11000000101001100000100100011001;
assign x[2142]= 32'b11000000101010100000100100110010;
assign x[2143]= 32'b11000000101011100000100101001011;
assign x[2144]= 32'b11000000101100010000100101100100;
assign x[2145]= 32'b11000000101101010000100101111100;
assign x[2146]= 32'b11000000101110010000100110010101;
assign x[2147]= 32'b11000000101111010000100110101110;
assign x[2148]= 32'b11000000110000000000100111000111;
assign x[2149]= 32'b11000000110001000000100111100000;
assign x[2150]= 32'b11000000110010000000100111111001;
assign x[2151]= 32'b11000000110011000000101000010001;
assign x[2152]= 32'b11000000110100000000101000101010;
assign x[2153]= 32'b11000000110101000000101001000011;
assign x[2154]= 32'b11000000110110000000101001011100;
assign x[2155]= 32'b11000000110111000000101001110101;
assign x[2156]= 32'b11000000111000000000101010001101;
assign x[2157]= 32'b11000000111001000000101010100110;
assign x[2158]= 32'b11000000111010010000101010111111;
assign x[2159]= 32'b11000000111011010000101011011000;
assign x[2160]= 32'b11000000111100010000101011110001;
assign x[2161]= 32'b11000000111101100000101100001001;
assign x[2162]= 32'b11000000111110100000101100100010;
assign x[2163]= 32'b11000000111111100000101100111011;
assign x[2164]= 32'b11000001000000110000101101010100;
assign x[2165]= 32'b11000001000001110000101101101100;
assign x[2166]= 32'b11000001000011000000101110000101;
assign x[2167]= 32'b11000001000100000000101110011110;
assign x[2168]= 32'b11000001000101010000101110110110;
assign x[2169]= 32'b11000001000110010000101111001111;
assign x[2170]= 32'b11000001000111100000101111101000;
assign x[2171]= 32'b11000001001000110000110000000001;
assign x[2172]= 32'b11000001001010000000110000011001;
assign x[2173]= 32'b11000001001011000000110000110010;
assign x[2174]= 32'b11000001001100010000110001001011;
assign x[2175]= 32'b11000001001101100000110001100011;
assign x[2176]= 32'b11000001001110110000110001111100;
assign x[2177]= 32'b11000001010000000000110010010101;
assign x[2178]= 32'b11000001010001010000110010101101;
assign x[2179]= 32'b11000001010010100000110011000110;
assign x[2180]= 32'b11000001010011110000110011011110;
assign x[2181]= 32'b11000001010101000000110011110111;
assign x[2182]= 32'b11000001010110010000110100010000;
assign x[2183]= 32'b11000001010111100000110100101000;
assign x[2184]= 32'b11000001011000110000110101000001;
assign x[2185]= 32'b11000001011010000000110101011001;
assign x[2186]= 32'b11000001011011100000110101110010;
assign x[2187]= 32'b11000001011100110000110110001011;
assign x[2188]= 32'b11000001011110000000110110100011;
assign x[2189]= 32'b11000001011111100000110110111100;
assign x[2190]= 32'b11000001100000110000110111010100;
assign x[2191]= 32'b11000001100010010000110111101101;
assign x[2192]= 32'b11000001100011100000111000000101;
assign x[2193]= 32'b11000001100101000000111000011110;
assign x[2194]= 32'b11000001100110010000111000110110;
assign x[2195]= 32'b11000001100111110000111001001111;
assign x[2196]= 32'b11000001101001000000111001100111;
assign x[2197]= 32'b11000001101010100000111010000000;
assign x[2198]= 32'b11000001101100000000111010011000;
assign x[2199]= 32'b11000001101101100000111010110001;
assign x[2200]= 32'b11000001101110110000111011001001;
assign x[2201]= 32'b11000001110000010000111011100010;
assign x[2202]= 32'b11000001110001110000111011111010;
assign x[2203]= 32'b11000001110011010000111100010010;
assign x[2204]= 32'b11000001110100110000111100101011;
assign x[2205]= 32'b11000001110110010000111101000011;
assign x[2206]= 32'b11000001110111110000111101011100;
assign x[2207]= 32'b11000001111001010000111101110100;
assign x[2208]= 32'b11000001111010110000111110001100;
assign x[2209]= 32'b11000001111100010000111110100101;
assign x[2210]= 32'b11000001111101110000111110111101;
assign x[2211]= 32'b11000001111111010000111111010110;
assign x[2212]= 32'b11000010000001000000111111101110;
assign x[2213]= 32'b11000010000010100001000000000110;
assign x[2214]= 32'b11000010000100000001000000011111;
assign x[2215]= 32'b11000010000101110001000000110111;
assign x[2216]= 32'b11000010000111010001000001001111;
assign x[2217]= 32'b11000010001000110001000001101000;
assign x[2218]= 32'b11000010001010100001000010000000;
assign x[2219]= 32'b11000010001100000001000010011000;
assign x[2220]= 32'b11000010001101110001000010110000;
assign x[2221]= 32'b11000010001111100001000011001001;
assign x[2222]= 32'b11000010010001000001000011100001;
assign x[2223]= 32'b11000010010010110001000011111001;
assign x[2224]= 32'b11000010010100010001000100010001;
assign x[2225]= 32'b11000010010110000001000100101010;
assign x[2226]= 32'b11000010010111110001000101000010;
assign x[2227]= 32'b11000010011001100001000101011010;
assign x[2228]= 32'b11000010011011010001000101110010;
assign x[2229]= 32'b11000010011100110001000110001010;
assign x[2230]= 32'b11000010011110100001000110100010;
assign x[2231]= 32'b11000010100000010001000110111011;
assign x[2232]= 32'b11000010100010000001000111010011;
assign x[2233]= 32'b11000010100011110001000111101011;
assign x[2234]= 32'b11000010100101100001001000000011;
assign x[2235]= 32'b11000010100111010001001000011011;
assign x[2236]= 32'b11000010101001010001001000110011;
assign x[2237]= 32'b11000010101011000001001001001011;
assign x[2238]= 32'b11000010101100110001001001100011;
assign x[2239]= 32'b11000010101110100001001001111011;
assign x[2240]= 32'b11000010110000010001001010010100;
assign x[2241]= 32'b11000010110010010001001010101100;
assign x[2242]= 32'b11000010110100000001001011000100;
assign x[2243]= 32'b11000010110110000001001011011100;
assign x[2244]= 32'b11000010110111110001001011110100;
assign x[2245]= 32'b11000010111001100001001100001100;
assign x[2246]= 32'b11000010111011100001001100100100;
assign x[2247]= 32'b11000010111101010001001100111100;
assign x[2248]= 32'b11000010111111010001001101010100;
assign x[2249]= 32'b11000011000001010001001101101100;
assign x[2250]= 32'b11000011000011000001001110000011;
assign x[2251]= 32'b11000011000101000001001110011011;
assign x[2252]= 32'b11000011000111000001001110110011;
assign x[2253]= 32'b11000011001000110001001111001011;
assign x[2254]= 32'b11000011001010110001001111100011;
assign x[2255]= 32'b11000011001100110001001111111011;
assign x[2256]= 32'b11000011001110110001010000010011;
assign x[2257]= 32'b11000011010000110001010000101011;
assign x[2258]= 32'b11000011010010110001010001000011;
assign x[2259]= 32'b11000011010100110001010001011010;
assign x[2260]= 32'b11000011010110110001010001110010;
assign x[2261]= 32'b11000011011000110001010010001010;
assign x[2262]= 32'b11000011011010110001010010100010;
assign x[2263]= 32'b11000011011100110001010010111010;
assign x[2264]= 32'b11000011011110110001010011010001;
assign x[2265]= 32'b11000011100000110001010011101001;
assign x[2266]= 32'b11000011100011000001010100000001;
assign x[2267]= 32'b11000011100101000001010100011001;
assign x[2268]= 32'b11000011100111000001010100110000;
assign x[2269]= 32'b11000011101001010001010101001000;
assign x[2270]= 32'b11000011101011010001010101100000;
assign x[2271]= 32'b11000011101101010001010101110111;
assign x[2272]= 32'b11000011101111100001010110001111;
assign x[2273]= 32'b11000011110001100001010110100111;
assign x[2274]= 32'b11000011110011110001010110111110;
assign x[2275]= 32'b11000011110101110001010111010110;
assign x[2276]= 32'b11000011111000000001010111101110;
assign x[2277]= 32'b11000011111010010001011000000101;
assign x[2278]= 32'b11000011111100010001011000011101;
assign x[2279]= 32'b11000011111110100001011000110100;
assign x[2280]= 32'b11000100000000110001011001001100;
assign x[2281]= 32'b11000100000010110001011001100100;
assign x[2282]= 32'b11000100000101000001011001111011;
assign x[2283]= 32'b11000100000111010001011010010011;
assign x[2284]= 32'b11000100001001100001011010101010;
assign x[2285]= 32'b11000100001011110001011011000010;
assign x[2286]= 32'b11000100001110000001011011011001;
assign x[2287]= 32'b11000100010000010001011011110001;
assign x[2288]= 32'b11000100010010100001011100001000;
assign x[2289]= 32'b11000100010100110001011100011111;
assign x[2290]= 32'b11000100010111000001011100110111;
assign x[2291]= 32'b11000100011001010001011101001110;
assign x[2292]= 32'b11000100011011100001011101100110;
assign x[2293]= 32'b11000100011110000001011101111101;
assign x[2294]= 32'b11000100100000010001011110010100;
assign x[2295]= 32'b11000100100010100001011110101100;
assign x[2296]= 32'b11000100100100110001011111000011;
assign x[2297]= 32'b11000100100111010001011111011010;
assign x[2298]= 32'b11000100101001100001011111110010;
assign x[2299]= 32'b11000100101100000001100000001001;
assign x[2300]= 32'b11000100101110010001100000100000;
assign x[2301]= 32'b11000100110000100001100000111000;
assign x[2302]= 32'b11000100110011000001100001001111;
assign x[2303]= 32'b11000100110101100001100001100110;
assign x[2304]= 32'b11000100110111110001100001111101;
assign x[2305]= 32'b11000100111010010001100010010101;
assign x[2306]= 32'b11000100111100100001100010101100;
assign x[2307]= 32'b11000100111111000001100011000011;
assign x[2308]= 32'b11000101000001100001100011011010;
assign x[2309]= 32'b11000101000100000001100011110001;
assign x[2310]= 32'b11000101000110100001100100001000;
assign x[2311]= 32'b11000101001000110001100100100000;
assign x[2312]= 32'b11000101001011010001100100110111;
assign x[2313]= 32'b11000101001101110001100101001110;
assign x[2314]= 32'b11000101010000010001100101100101;
assign x[2315]= 32'b11000101010010110001100101111100;
assign x[2316]= 32'b11000101010101010001100110010011;
assign x[2317]= 32'b11000101010111110001100110101010;
assign x[2318]= 32'b11000101011010010001100111000001;
assign x[2319]= 32'b11000101011100110001100111011000;
assign x[2320]= 32'b11000101011111100001100111101111;
assign x[2321]= 32'b11000101100010000001101000000110;
assign x[2322]= 32'b11000101100100100001101000011101;
assign x[2323]= 32'b11000101100111000001101000110100;
assign x[2324]= 32'b11000101101001110001101001001011;
assign x[2325]= 32'b11000101101100010001101001100010;
assign x[2326]= 32'b11000101101110110001101001111001;
assign x[2327]= 32'b11000101110001100001101010001111;
assign x[2328]= 32'b11000101110100000001101010100110;
assign x[2329]= 32'b11000101110110110001101010111101;
assign x[2330]= 32'b11000101111001010001101011010100;
assign x[2331]= 32'b11000101111100000001101011101011;
assign x[2332]= 32'b11000101111110100001101100000010;
assign x[2333]= 32'b11000110000001010001101100011000;
assign x[2334]= 32'b11000110000100000001101100101111;
assign x[2335]= 32'b11000110000110100001101101000110;
assign x[2336]= 32'b11000110001001010001101101011101;
assign x[2337]= 32'b11000110001100000001101101110011;
assign x[2338]= 32'b11000110001110110001101110001010;
assign x[2339]= 32'b11000110010001010001101110100001;
assign x[2340]= 32'b11000110010100000001101110110111;
assign x[2341]= 32'b11000110010110110001101111001110;
assign x[2342]= 32'b11000110011001100001101111100101;
assign x[2343]= 32'b11000110011100010001101111111011;
assign x[2344]= 32'b11000110011111000001110000010010;
assign x[2345]= 32'b11000110100001110001110000101000;
assign x[2346]= 32'b11000110100100100001110000111111;
assign x[2347]= 32'b11000110100111010001110001010101;
assign x[2348]= 32'b11000110101010000001110001101100;
assign x[2349]= 32'b11000110101101000001110010000011;
assign x[2350]= 32'b11000110101111110001110010011001;
assign x[2351]= 32'b11000110110010100001110010101111;
assign x[2352]= 32'b11000110110101010001110011000110;
assign x[2353]= 32'b11000110111000010001110011011100;
assign x[2354]= 32'b11000110111011000001110011110011;
assign x[2355]= 32'b11000110111101110001110100001001;
assign x[2356]= 32'b11000111000000110001110100100000;
assign x[2357]= 32'b11000111000011100001110100110110;
assign x[2358]= 32'b11000111000110100001110101001100;
assign x[2359]= 32'b11000111001001010001110101100011;
assign x[2360]= 32'b11000111001100010001110101111001;
assign x[2361]= 32'b11000111001111010001110110001111;
assign x[2362]= 32'b11000111010010000001110110100110;
assign x[2363]= 32'b11000111010101000001110110111100;
assign x[2364]= 32'b11000111010111110001110111010010;
assign x[2365]= 32'b11000111011010110001110111101000;
assign x[2366]= 32'b11000111011101110001110111111110;
assign x[2367]= 32'b11000111100000110001111000010101;
assign x[2368]= 32'b11000111100011110001111000101011;
assign x[2369]= 32'b11000111100110100001111001000001;
assign x[2370]= 32'b11000111101001100001111001010111;
assign x[2371]= 32'b11000111101100100001111001101101;
assign x[2372]= 32'b11000111101111100001111010000011;
assign x[2373]= 32'b11000111110010100001111010011001;
assign x[2374]= 32'b11000111110101100001111010110000;
assign x[2375]= 32'b11000111111000100001111011000110;
assign x[2376]= 32'b11000111111011100001111011011100;
assign x[2377]= 32'b11000111111110110001111011110010;
assign x[2378]= 32'b11001000000001110001111100001000;
assign x[2379]= 32'b11001000000100110001111100011110;
assign x[2380]= 32'b11001000000111110001111100110100;
assign x[2381]= 32'b11001000001010110001111101001001;
assign x[2382]= 32'b11001000001110000001111101011111;
assign x[2383]= 32'b11001000010001000001111101110101;
assign x[2384]= 32'b11001000010100000001111110001011;
assign x[2385]= 32'b11001000010111010001111110100001;
assign x[2386]= 32'b11001000011010010001111110110111;
assign x[2387]= 32'b11001000011101100001111111001101;
assign x[2388]= 32'b11001000100000100001111111100010;
assign x[2389]= 32'b11001000100011110001111111111000;
assign x[2390]= 32'b11001000100110110010000000001110;
assign x[2391]= 32'b11001000101010000010000000100100;
assign x[2392]= 32'b11001000101101010010000000111001;
assign x[2393]= 32'b11001000110000010010000001001111;
assign x[2394]= 32'b11001000110011100010000001100101;
assign x[2395]= 32'b11001000110110110010000001111011;
assign x[2396]= 32'b11001000111010000010000010010000;
assign x[2397]= 32'b11001000111101000010000010100110;
assign x[2398]= 32'b11001001000000010010000010111011;
assign x[2399]= 32'b11001001000011100010000011010001;
assign x[2400]= 32'b11001001000110110010000011100111;
assign x[2401]= 32'b11001001001010000010000011111100;
assign x[2402]= 32'b11001001001101010010000100010010;
assign x[2403]= 32'b11001001010000100010000100100111;
assign x[2404]= 32'b11001001010011110010000100111101;
assign x[2405]= 32'b11001001010111000010000101010010;
assign x[2406]= 32'b11001001011010010010000101101000;
assign x[2407]= 32'b11001001011101100010000101111101;
assign x[2408]= 32'b11001001100000110010000110010010;
assign x[2409]= 32'b11001001100100010010000110101000;
assign x[2410]= 32'b11001001100111100010000110111101;
assign x[2411]= 32'b11001001101010110010000111010010;
assign x[2412]= 32'b11001001101110000010000111101000;
assign x[2413]= 32'b11001001110001100010000111111101;
assign x[2414]= 32'b11001001110100110010001000010010;
assign x[2415]= 32'b11001001111000000010001000101000;
assign x[2416]= 32'b11001001111011100010001000111101;
assign x[2417]= 32'b11001001111110110010001001010010;
assign x[2418]= 32'b11001010000010010010001001100111;
assign x[2419]= 32'b11001010000101100010001001111101;
assign x[2420]= 32'b11001010001001000010001010010010;
assign x[2421]= 32'b11001010001100100010001010100111;
assign x[2422]= 32'b11001010001111110010001010111100;
assign x[2423]= 32'b11001010010011010010001011010001;
assign x[2424]= 32'b11001010010110110010001011100110;
assign x[2425]= 32'b11001010011010000010001011111011;
assign x[2426]= 32'b11001010011101100010001100010000;
assign x[2427]= 32'b11001010100001000010001100100101;
assign x[2428]= 32'b11001010100100100010001100111010;
assign x[2429]= 32'b11001010100111110010001101001111;
assign x[2430]= 32'b11001010101011010010001101100100;
assign x[2431]= 32'b11001010101110110010001101111001;
assign x[2432]= 32'b11001010110010010010001110001110;
assign x[2433]= 32'b11001010110101110010001110100011;
assign x[2434]= 32'b11001010111001010010001110111000;
assign x[2435]= 32'b11001010111100110010001111001101;
assign x[2436]= 32'b11001011000000010010001111100001;
assign x[2437]= 32'b11001011000011110010001111110110;
assign x[2438]= 32'b11001011000111100010010000001011;
assign x[2439]= 32'b11001011001011000010010000100000;
assign x[2440]= 32'b11001011001110100010010000110100;
assign x[2441]= 32'b11001011010010000010010001001001;
assign x[2442]= 32'b11001011010101100010010001011110;
assign x[2443]= 32'b11001011011001010010010001110011;
assign x[2444]= 32'b11001011011100110010010010000111;
assign x[2445]= 32'b11001011100000010010010010011100;
assign x[2446]= 32'b11001011100100000010010010110000;
assign x[2447]= 32'b11001011100111100010010011000101;
assign x[2448]= 32'b11001011101011010010010011011010;
assign x[2449]= 32'b11001011101110110010010011101110;
assign x[2450]= 32'b11001011110010100010010100000011;
assign x[2451]= 32'b11001011110110000010010100010111;
assign x[2452]= 32'b11001011111001110010010100101100;
assign x[2453]= 32'b11001011111101010010010101000000;
assign x[2454]= 32'b11001100000001000010010101010100;
assign x[2455]= 32'b11001100000100110010010101101001;
assign x[2456]= 32'b11001100001000010010010101111101;
assign x[2457]= 32'b11001100001100000010010110010010;
assign x[2458]= 32'b11001100001111110010010110100110;
assign x[2459]= 32'b11001100010011100010010110111010;
assign x[2460]= 32'b11001100010111010010010111001111;
assign x[2461]= 32'b11001100011010110010010111100011;
assign x[2462]= 32'b11001100011110100010010111110111;
assign x[2463]= 32'b11001100100010010010011000001011;
assign x[2464]= 32'b11001100100110000010011000011111;
assign x[2465]= 32'b11001100101001110010011000110100;
assign x[2466]= 32'b11001100101101100010011001001000;
assign x[2467]= 32'b11001100110001010010011001011100;
assign x[2468]= 32'b11001100110101000010011001110000;
assign x[2469]= 32'b11001100111000110010011010000100;
assign x[2470]= 32'b11001100111100110010011010011000;
assign x[2471]= 32'b11001101000000100010011010101100;
assign x[2472]= 32'b11001101000100010010011011000000;
assign x[2473]= 32'b11001101001000000010011011010100;
assign x[2474]= 32'b11001101001100000010011011101000;
assign x[2475]= 32'b11001101001111110010011011111100;
assign x[2476]= 32'b11001101010011100010011100010000;
assign x[2477]= 32'b11001101010111010010011100100100;
assign x[2478]= 32'b11001101011011010010011100111000;
assign x[2479]= 32'b11001101011111000010011101001100;
assign x[2480]= 32'b11001101100011000010011101011111;
assign x[2481]= 32'b11001101100110110010011101110011;
assign x[2482]= 32'b11001101101010110010011110000111;
assign x[2483]= 32'b11001101101110100010011110011011;
assign x[2484]= 32'b11001101110010100010011110101111;
assign x[2485]= 32'b11001101110110010010011111000010;
assign x[2486]= 32'b11001101111010010010011111010110;
assign x[2487]= 32'b11001101111110010010011111101010;
assign x[2488]= 32'b11001110000010000010011111111101;
assign x[2489]= 32'b11001110000110000010100000010001;
assign x[2490]= 32'b11001110001010000010100000100100;
assign x[2491]= 32'b11001110001110000010100000111000;
assign x[2492]= 32'b11001110010001110010100001001011;
assign x[2493]= 32'b11001110010101110010100001011111;
assign x[2494]= 32'b11001110011001110010100001110010;
assign x[2495]= 32'b11001110011101110010100010000110;
assign x[2496]= 32'b11001110100001110010100010011001;
assign x[2497]= 32'b11001110100101110010100010101101;
assign x[2498]= 32'b11001110101001110010100011000000;
assign x[2499]= 32'b11001110101101110010100011010100;
assign x[2500]= 32'b11001110110001110010100011100111;
assign x[2501]= 32'b11001110110101110010100011111010;
assign x[2502]= 32'b11001110111001110010100100001110;
assign x[2503]= 32'b11001110111101110010100100100001;
assign x[2504]= 32'b11001111000001110010100100110100;
assign x[2505]= 32'b11001111000110000010100101000111;
assign x[2506]= 32'b11001111001010000010100101011010;
assign x[2507]= 32'b11001111001110000010100101101110;
assign x[2508]= 32'b11001111010010000010100110000001;
assign x[2509]= 32'b11001111010110010010100110010100;
assign x[2510]= 32'b11001111011010010010100110100111;
assign x[2511]= 32'b11001111011110010010100110111010;
assign x[2512]= 32'b11001111100010100010100111001101;
assign x[2513]= 32'b11001111100110100010100111100000;
assign x[2514]= 32'b11001111101010110010100111110011;
assign x[2515]= 32'b11001111101110110010101000000110;
assign x[2516]= 32'b11001111110011000010101000011001;
assign x[2517]= 32'b11001111110111000010101000101100;
assign x[2518]= 32'b11001111111011010010101000111111;
assign x[2519]= 32'b11001111111111100010101001010010;
assign x[2520]= 32'b11010000000011100010101001100101;
assign x[2521]= 32'b11010000000111110010101001110111;
assign x[2522]= 32'b11010000001100000010101010001010;
assign x[2523]= 32'b11010000010000000010101010011101;
assign x[2524]= 32'b11010000010100010010101010110000;
assign x[2525]= 32'b11010000011000100010101011000010;
assign x[2526]= 32'b11010000011100110010101011010101;
assign x[2527]= 32'b11010000100000110010101011101000;
assign x[2528]= 32'b11010000100101000010101011111010;
assign x[2529]= 32'b11010000101001010010101100001101;
assign x[2530]= 32'b11010000101101100010101100100000;
assign x[2531]= 32'b11010000110001110010101100110010;
assign x[2532]= 32'b11010000110110000010101101000101;
assign x[2533]= 32'b11010000111010010010101101010111;
assign x[2534]= 32'b11010000111110100010101101101010;
assign x[2535]= 32'b11010001000010110010101101111100;
assign x[2536]= 32'b11010001000111000010101110001110;
assign x[2537]= 32'b11010001001011010010101110100001;
assign x[2538]= 32'b11010001001111100010101110110011;
assign x[2539]= 32'b11010001010100000010101111000110;
assign x[2540]= 32'b11010001011000010010101111011000;
assign x[2541]= 32'b11010001011100100010101111101010;
assign x[2542]= 32'b11010001100000110010101111111100;
assign x[2543]= 32'b11010001100101010010110000001111;
assign x[2544]= 32'b11010001101001100010110000100001;
assign x[2545]= 32'b11010001101101110010110000110011;
assign x[2546]= 32'b11010001110010010010110001000101;
assign x[2547]= 32'b11010001110110100010110001010111;
assign x[2548]= 32'b11010001111010110010110001101010;
assign x[2549]= 32'b11010001111111010010110001111100;
assign x[2550]= 32'b11010010000011100010110010001110;
assign x[2551]= 32'b11010010001000000010110010100000;
assign x[2552]= 32'b11010010001100010010110010110010;
assign x[2553]= 32'b11010010010000110010110011000100;
assign x[2554]= 32'b11010010010101010010110011010110;
assign x[2555]= 32'b11010010011001100010110011101000;
assign x[2556]= 32'b11010010011110000010110011111001;
assign x[2557]= 32'b11010010100010100010110100001011;
assign x[2558]= 32'b11010010100110110010110100011101;
assign x[2559]= 32'b11010010101011010010110100101111;
assign x[2560]= 32'b11010010101111110010110101000001;
assign x[2561]= 32'b11010010110100010010110101010010;
assign x[2562]= 32'b11010010111000100010110101100100;
assign x[2563]= 32'b11010010111101000010110101110110;
assign x[2564]= 32'b11010011000001100010110110001000;
assign x[2565]= 32'b11010011000110000010110110011001;
assign x[2566]= 32'b11010011001010100010110110101011;
assign x[2567]= 32'b11010011001111000010110110111100;
assign x[2568]= 32'b11010011010011100010110111001110;
assign x[2569]= 32'b11010011011000000010110111100000;
assign x[2570]= 32'b11010011011100100010110111110001;
assign x[2571]= 32'b11010011100001000010111000000011;
assign x[2572]= 32'b11010011100101100010111000010100;
assign x[2573]= 32'b11010011101010000010111000100101;
assign x[2574]= 32'b11010011101110100010111000110111;
assign x[2575]= 32'b11010011110011000010111001001000;
assign x[2576]= 32'b11010011110111110010111001011010;
assign x[2577]= 32'b11010011111100010010111001101011;
assign x[2578]= 32'b11010100000000110010111001111100;
assign x[2579]= 32'b11010100000101010010111010001101;
assign x[2580]= 32'b11010100001010000010111010011111;
assign x[2581]= 32'b11010100001110100010111010110000;
assign x[2582]= 32'b11010100010011000010111011000001;
assign x[2583]= 32'b11010100010111110010111011010010;
assign x[2584]= 32'b11010100011100010010111011100011;
assign x[2585]= 32'b11010100100000110010111011110100;
assign x[2586]= 32'b11010100100101100010111100000101;
assign x[2587]= 32'b11010100101010000010111100010110;
assign x[2588]= 32'b11010100101110110010111100101000;
assign x[2589]= 32'b11010100110011010010111100111000;
assign x[2590]= 32'b11010100111000000010111101001001;
assign x[2591]= 32'b11010100111100110010111101011010;
assign x[2592]= 32'b11010101000001010010111101101011;
assign x[2593]= 32'b11010101000110000010111101111100;
assign x[2594]= 32'b11010101001010100010111110001101;
assign x[2595]= 32'b11010101001111010010111110011110;
assign x[2596]= 32'b11010101010100000010111110101111;
assign x[2597]= 32'b11010101011000110010111110111111;
assign x[2598]= 32'b11010101011101010010111111010000;
assign x[2599]= 32'b11010101100010000010111111100001;
assign x[2600]= 32'b11010101100110110010111111110001;
assign x[2601]= 32'b11010101101011100011000000000010;
assign x[2602]= 32'b11010101110000010011000000010011;
assign x[2603]= 32'b11010101110101000011000000100011;
assign x[2604]= 32'b11010101111001100011000000110100;
assign x[2605]= 32'b11010101111110010011000001000100;
assign x[2606]= 32'b11010110000011000011000001010101;
assign x[2607]= 32'b11010110000111110011000001100101;
assign x[2608]= 32'b11010110001100100011000001110110;
assign x[2609]= 32'b11010110010001010011000010000110;
assign x[2610]= 32'b11010110010110010011000010010110;
assign x[2611]= 32'b11010110011011000011000010100111;
assign x[2612]= 32'b11010110011111110011000010110111;
assign x[2613]= 32'b11010110100100100011000011000111;
assign x[2614]= 32'b11010110101001010011000011011000;
assign x[2615]= 32'b11010110101110000011000011101000;
assign x[2616]= 32'b11010110110010110011000011111000;
assign x[2617]= 32'b11010110110111110011000100001000;
assign x[2618]= 32'b11010110111100100011000100011000;
assign x[2619]= 32'b11010111000001010011000100101000;
assign x[2620]= 32'b11010111000110010011000100111000;
assign x[2621]= 32'b11010111001011000011000101001001;
assign x[2622]= 32'b11010111001111110011000101011001;
assign x[2623]= 32'b11010111010100110011000101101001;
assign x[2624]= 32'b11010111011001100011000101111001;
assign x[2625]= 32'b11010111011110100011000110001000;
assign x[2626]= 32'b11010111100011010011000110011000;
assign x[2627]= 32'b11010111101000000011000110101000;
assign x[2628]= 32'b11010111101101000011000110111000;
assign x[2629]= 32'b11010111110010000011000111001000;
assign x[2630]= 32'b11010111110110110011000111011000;
assign x[2631]= 32'b11010111111011110011000111100111;
assign x[2632]= 32'b11011000000000100011000111110111;
assign x[2633]= 32'b11011000000101100011001000000111;
assign x[2634]= 32'b11011000001010100011001000010110;
assign x[2635]= 32'b11011000001111010011001000100110;
assign x[2636]= 32'b11011000010100010011001000110110;
assign x[2637]= 32'b11011000011001010011001001000101;
assign x[2638]= 32'b11011000011110000011001001010101;
assign x[2639]= 32'b11011000100011000011001001100100;
assign x[2640]= 32'b11011000101000000011001001110100;
assign x[2641]= 32'b11011000101101000011001010000011;
assign x[2642]= 32'b11011000110010000011001010010011;
assign x[2643]= 32'b11011000110111000011001010100010;
assign x[2644]= 32'b11011000111011110011001010110001;
assign x[2645]= 32'b11011001000000110011001011000001;
assign x[2646]= 32'b11011001000101110011001011010000;
assign x[2647]= 32'b11011001001010110011001011011111;
assign x[2648]= 32'b11011001001111110011001011101110;
assign x[2649]= 32'b11011001010100110011001011111110;
assign x[2650]= 32'b11011001011001110011001100001101;
assign x[2651]= 32'b11011001011110110011001100011100;
assign x[2652]= 32'b11011001100011110011001100101011;
assign x[2653]= 32'b11011001101001000011001100111010;
assign x[2654]= 32'b11011001101110000011001101001001;
assign x[2655]= 32'b11011001110011000011001101011000;
assign x[2656]= 32'b11011001111000000011001101100111;
assign x[2657]= 32'b11011001111101000011001101110110;
assign x[2658]= 32'b11011010000010000011001110000101;
assign x[2659]= 32'b11011010000111010011001110010100;
assign x[2660]= 32'b11011010001100010011001110100011;
assign x[2661]= 32'b11011010010001010011001110110010;
assign x[2662]= 32'b11011010010110100011001111000001;
assign x[2663]= 32'b11011010011011100011001111001111;
assign x[2664]= 32'b11011010100000100011001111011110;
assign x[2665]= 32'b11011010100101110011001111101101;
assign x[2666]= 32'b11011010101010110011001111111011;
assign x[2667]= 32'b11011010101111110011010000001010;
assign x[2668]= 32'b11011010110101000011010000011001;
assign x[2669]= 32'b11011010111010000011010000100111;
assign x[2670]= 32'b11011010111111010011010000110110;
assign x[2671]= 32'b11011011000100010011010001000100;
assign x[2672]= 32'b11011011001001100011010001010011;
assign x[2673]= 32'b11011011001110110011010001100001;
assign x[2674]= 32'b11011011010011110011010001110000;
assign x[2675]= 32'b11011011011001000011010001111110;
assign x[2676]= 32'b11011011011110000011010010001100;
assign x[2677]= 32'b11011011100011010011010010011011;
assign x[2678]= 32'b11011011101000100011010010101001;
assign x[2679]= 32'b11011011101101100011010010110111;
assign x[2680]= 32'b11011011110010110011010011000110;
assign x[2681]= 32'b11011011111000000011010011010100;
assign x[2682]= 32'b11011011111101010011010011100010;
assign x[2683]= 32'b11011100000010010011010011110000;
assign x[2684]= 32'b11011100000111100011010011111110;
assign x[2685]= 32'b11011100001100110011010100001100;
assign x[2686]= 32'b11011100010010000011010100011010;
assign x[2687]= 32'b11011100010111010011010100101000;
assign x[2688]= 32'b11011100011100100011010100110110;
assign x[2689]= 32'b11011100100001100011010101000100;
assign x[2690]= 32'b11011100100110110011010101010010;
assign x[2691]= 32'b11011100101100000011010101100000;
assign x[2692]= 32'b11011100110001010011010101101110;
assign x[2693]= 32'b11011100110110100011010101111100;
assign x[2694]= 32'b11011100111011110011010110001001;
assign x[2695]= 32'b11011101000001000011010110010111;
assign x[2696]= 32'b11011101000110010011010110100101;
assign x[2697]= 32'b11011101001011100011010110110011;
assign x[2698]= 32'b11011101010001000011010111000000;
assign x[2699]= 32'b11011101010110010011010111001110;
assign x[2700]= 32'b11011101011011100011010111011100;
assign x[2701]= 32'b11011101100000110011010111101001;
assign x[2702]= 32'b11011101100110000011010111110111;
assign x[2703]= 32'b11011101101011010011011000000100;
assign x[2704]= 32'b11011101110000110011011000010010;
assign x[2705]= 32'b11011101110110000011011000011111;
assign x[2706]= 32'b11011101111011010011011000101100;
assign x[2707]= 32'b11011110000000100011011000111010;
assign x[2708]= 32'b11011110000110000011011001000111;
assign x[2709]= 32'b11011110001011010011011001010100;
assign x[2710]= 32'b11011110010000100011011001100010;
assign x[2711]= 32'b11011110010110000011011001101111;
assign x[2712]= 32'b11011110011011010011011001111100;
assign x[2713]= 32'b11011110100000110011011010001001;
assign x[2714]= 32'b11011110100110000011011010010110;
assign x[2715]= 32'b11011110101011010011011010100100;
assign x[2716]= 32'b11011110110000110011011010110001;
assign x[2717]= 32'b11011110110110000011011010111110;
assign x[2718]= 32'b11011110111011100011011011001011;
assign x[2719]= 32'b11011111000000110011011011011000;
assign x[2720]= 32'b11011111000110010011011011100101;
assign x[2721]= 32'b11011111001011110011011011110001;
assign x[2722]= 32'b11011111010001000011011011111110;
assign x[2723]= 32'b11011111010110100011011100001011;
assign x[2724]= 32'b11011111011011110011011100011000;
assign x[2725]= 32'b11011111100001010011011100100101;
assign x[2726]= 32'b11011111100110110011011100110001;
assign x[2727]= 32'b11011111101100000011011100111110;
assign x[2728]= 32'b11011111110001100011011101001011;
assign x[2729]= 32'b11011111110111000011011101010111;
assign x[2730]= 32'b11011111111100010011011101100100;
assign x[2731]= 32'b11100000000001110011011101110001;
assign x[2732]= 32'b11100000000111010011011101111101;
assign x[2733]= 32'b11100000001100110011011110001010;
assign x[2734]= 32'b11100000010010010011011110010110;
assign x[2735]= 32'b11100000010111100011011110100011;
assign x[2736]= 32'b11100000011101000011011110101111;
assign x[2737]= 32'b11100000100010100011011110111011;
assign x[2738]= 32'b11100000101000000011011111001000;
assign x[2739]= 32'b11100000101101100011011111010100;
assign x[2740]= 32'b11100000110011000011011111100000;
assign x[2741]= 32'b11100000111000100011011111101101;
assign x[2742]= 32'b11100000111110000011011111111001;
assign x[2743]= 32'b11100001000011100011100000000101;
assign x[2744]= 32'b11100001001001000011100000010001;
assign x[2745]= 32'b11100001001110100011100000011101;
assign x[2746]= 32'b11100001010100000011100000101001;
assign x[2747]= 32'b11100001011001100011100000110101;
assign x[2748]= 32'b11100001011111000011100001000001;
assign x[2749]= 32'b11100001100100100011100001001101;
assign x[2750]= 32'b11100001101010000011100001011001;
assign x[2751]= 32'b11100001101111100011100001100101;
assign x[2752]= 32'b11100001110101010011100001110001;
assign x[2753]= 32'b11100001111010110011100001111101;
assign x[2754]= 32'b11100010000000010011100010001001;
assign x[2755]= 32'b11100010000101110011100010010100;
assign x[2756]= 32'b11100010001011010011100010100000;
assign x[2757]= 32'b11100010010001000011100010101100;
assign x[2758]= 32'b11100010010110100011100010110111;
assign x[2759]= 32'b11100010011100000011100011000011;
assign x[2760]= 32'b11100010100001110011100011001111;
assign x[2761]= 32'b11100010100111010011100011011010;
assign x[2762]= 32'b11100010101100110011100011100110;
assign x[2763]= 32'b11100010110010100011100011110001;
assign x[2764]= 32'b11100010111000000011100011111101;
assign x[2765]= 32'b11100010111101100011100100001000;
assign x[2766]= 32'b11100011000011010011100100010011;
assign x[2767]= 32'b11100011001000110011100100011111;
assign x[2768]= 32'b11100011001110100011100100101010;
assign x[2769]= 32'b11100011010100000011100100110101;
assign x[2770]= 32'b11100011011001110011100101000001;
assign x[2771]= 32'b11100011011111010011100101001100;
assign x[2772]= 32'b11100011100101000011100101010111;
assign x[2773]= 32'b11100011101010100011100101100010;
assign x[2774]= 32'b11100011110000010011100101101101;
assign x[2775]= 32'b11100011110101110011100101111000;
assign x[2776]= 32'b11100011111011100011100110000011;
assign x[2777]= 32'b11100100000001000011100110001110;
assign x[2778]= 32'b11100100000110110011100110011001;
assign x[2779]= 32'b11100100001100100011100110100100;
assign x[2780]= 32'b11100100010010000011100110101111;
assign x[2781]= 32'b11100100010111110011100110111010;
assign x[2782]= 32'b11100100011101100011100111000101;
assign x[2783]= 32'b11100100100011000011100111010000;
assign x[2784]= 32'b11100100101000110011100111011010;
assign x[2785]= 32'b11100100101110100011100111100101;
assign x[2786]= 32'b11100100110100000011100111110000;
assign x[2787]= 32'b11100100111001110011100111111011;
assign x[2788]= 32'b11100100111111100011101000000101;
assign x[2789]= 32'b11100101000101010011101000010000;
assign x[2790]= 32'b11100101001011000011101000011010;
assign x[2791]= 32'b11100101010000100011101000100101;
assign x[2792]= 32'b11100101010110010011101000101111;
assign x[2793]= 32'b11100101011100000011101000111010;
assign x[2794]= 32'b11100101100001110011101001000100;
assign x[2795]= 32'b11100101100111100011101001001111;
assign x[2796]= 32'b11100101101101010011101001011001;
assign x[2797]= 32'b11100101110011000011101001100011;
assign x[2798]= 32'b11100101111000110011101001101101;
assign x[2799]= 32'b11100101111110100011101001111000;
assign x[2800]= 32'b11100110000100010011101010000010;
assign x[2801]= 32'b11100110001010000011101010001100;
assign x[2802]= 32'b11100110001111110011101010010110;
assign x[2803]= 32'b11100110010101100011101010100000;
assign x[2804]= 32'b11100110011011010011101010101010;
assign x[2805]= 32'b11100110100001000011101010110100;
assign x[2806]= 32'b11100110100110110011101010111110;
assign x[2807]= 32'b11100110101100100011101011001000;
assign x[2808]= 32'b11100110110010010011101011010010;
assign x[2809]= 32'b11100110111000000011101011011100;
assign x[2810]= 32'b11100110111101110011101011100110;
assign x[2811]= 32'b11100111000011100011101011110000;
assign x[2812]= 32'b11100111001001010011101011111010;
assign x[2813]= 32'b11100111001111010011101100000011;
assign x[2814]= 32'b11100111010101000011101100001101;
assign x[2815]= 32'b11100111011010110011101100010111;
assign x[2816]= 32'b11100111100000100011101100100000;
assign x[2817]= 32'b11100111100110010011101100101010;
assign x[2818]= 32'b11100111101100010011101100110100;
assign x[2819]= 32'b11100111110010000011101100111101;
assign x[2820]= 32'b11100111110111110011101101000111;
assign x[2821]= 32'b11100111111101100011101101010000;
assign x[2822]= 32'b11101000000011100011101101011001;
assign x[2823]= 32'b11101000001001010011101101100011;
assign x[2824]= 32'b11101000001111000011101101101100;
assign x[2825]= 32'b11101000010101000011101101110101;
assign x[2826]= 32'b11101000011010110011101101111111;
assign x[2827]= 32'b11101000100000100011101110001000;
assign x[2828]= 32'b11101000100110100011101110010001;
assign x[2829]= 32'b11101000101100010011101110011010;
assign x[2830]= 32'b11101000110010010011101110100011;
assign x[2831]= 32'b11101000111000000011101110101101;
assign x[2832]= 32'b11101000111101110011101110110110;
assign x[2833]= 32'b11101001000011110011101110111111;
assign x[2834]= 32'b11101001001001100011101111001000;
assign x[2835]= 32'b11101001001111100011101111010001;
assign x[2836]= 32'b11101001010101010011101111011010;
assign x[2837]= 32'b11101001011011010011101111100010;
assign x[2838]= 32'b11101001100001000011101111101011;
assign x[2839]= 32'b11101001100111000011101111110100;
assign x[2840]= 32'b11101001101101000011101111111101;
assign x[2841]= 32'b11101001110010110011110000000110;
assign x[2842]= 32'b11101001111000110011110000001110;
assign x[2843]= 32'b11101001111110100011110000010111;
assign x[2844]= 32'b11101010000100100011110000100000;
assign x[2845]= 32'b11101010001010010011110000101000;
assign x[2846]= 32'b11101010010000010011110000110001;
assign x[2847]= 32'b11101010010110010011110000111001;
assign x[2848]= 32'b11101010011100000011110001000010;
assign x[2849]= 32'b11101010100010000011110001001010;
assign x[2850]= 32'b11101010101000000011110001010011;
assign x[2851]= 32'b11101010101101110011110001011011;
assign x[2852]= 32'b11101010110011110011110001100011;
assign x[2853]= 32'b11101010111001110011110001101100;
assign x[2854]= 32'b11101010111111110011110001110100;
assign x[2855]= 32'b11101011000101100011110001111100;
assign x[2856]= 32'b11101011001011100011110010000100;
assign x[2857]= 32'b11101011010001100011110010001100;
assign x[2858]= 32'b11101011010111100011110010010101;
assign x[2859]= 32'b11101011011101010011110010011101;
assign x[2860]= 32'b11101011100011010011110010100101;
assign x[2861]= 32'b11101011101001010011110010101101;
assign x[2862]= 32'b11101011101111010011110010110101;
assign x[2863]= 32'b11101011110101010011110010111101;
assign x[2864]= 32'b11101011111011010011110011000101;
assign x[2865]= 32'b11101100000001010011110011001100;
assign x[2866]= 32'b11101100000111000011110011010100;
assign x[2867]= 32'b11101100001101000011110011011100;
assign x[2868]= 32'b11101100010011000011110011100100;
assign x[2869]= 32'b11101100011001000011110011101100;
assign x[2870]= 32'b11101100011111000011110011110011;
assign x[2871]= 32'b11101100100101000011110011111011;
assign x[2872]= 32'b11101100101011000011110100000010;
assign x[2873]= 32'b11101100110001000011110100001010;
assign x[2874]= 32'b11101100110111000011110100010010;
assign x[2875]= 32'b11101100111101000011110100011001;
assign x[2876]= 32'b11101101000011000011110100100001;
assign x[2877]= 32'b11101101001001000011110100101000;
assign x[2878]= 32'b11101101001111000011110100101111;
assign x[2879]= 32'b11101101010101000011110100110111;
assign x[2880]= 32'b11101101011011000011110100111110;
assign x[2881]= 32'b11101101100001000011110101000101;
assign x[2882]= 32'b11101101100111000011110101001101;
assign x[2883]= 32'b11101101101101000011110101010100;
assign x[2884]= 32'b11101101110011000011110101011011;
assign x[2885]= 32'b11101101111001000011110101100010;
assign x[2886]= 32'b11101101111111000011110101101001;
assign x[2887]= 32'b11101110000101010011110101110000;
assign x[2888]= 32'b11101110001011010011110101110111;
assign x[2889]= 32'b11101110010001010011110101111110;
assign x[2890]= 32'b11101110010111010011110110000101;
assign x[2891]= 32'b11101110011101010011110110001100;
assign x[2892]= 32'b11101110100011010011110110010011;
assign x[2893]= 32'b11101110101001100011110110011010;
assign x[2894]= 32'b11101110101111100011110110100001;
assign x[2895]= 32'b11101110110101100011110110100111;
assign x[2896]= 32'b11101110111011100011110110101110;
assign x[2897]= 32'b11101111000001100011110110110101;
assign x[2898]= 32'b11101111000111110011110110111011;
assign x[2899]= 32'b11101111001101110011110111000010;
assign x[2900]= 32'b11101111010011110011110111001001;
assign x[2901]= 32'b11101111011001110011110111001111;
assign x[2902]= 32'b11101111100000000011110111010110;
assign x[2903]= 32'b11101111100110000011110111011100;
assign x[2904]= 32'b11101111101100000011110111100010;
assign x[2905]= 32'b11101111110010010011110111101001;
assign x[2906]= 32'b11101111111000010011110111101111;
assign x[2907]= 32'b11101111111110010011110111110101;
assign x[2908]= 32'b11110000000100100011110111111100;
assign x[2909]= 32'b11110000001010100011111000000010;
assign x[2910]= 32'b11110000010000100011111000001000;
assign x[2911]= 32'b11110000010110110011111000001110;
assign x[2912]= 32'b11110000011100110011111000010100;
assign x[2913]= 32'b11110000100010110011111000011011;
assign x[2914]= 32'b11110000101001000011111000100001;
assign x[2915]= 32'b11110000101111000011111000100111;
assign x[2916]= 32'b11110000110101010011111000101101;
assign x[2917]= 32'b11110000111011010011111000110011;
assign x[2918]= 32'b11110001000001010011111000111000;
assign x[2919]= 32'b11110001000111100011111000111110;
assign x[2920]= 32'b11110001001101100011111001000100;
assign x[2921]= 32'b11110001010011110011111001001010;
assign x[2922]= 32'b11110001011001110011111001010000;
assign x[2923]= 32'b11110001100000000011111001010101;
assign x[2924]= 32'b11110001100110000011111001011011;
assign x[2925]= 32'b11110001101100010011111001100001;
assign x[2926]= 32'b11110001110010010011111001100110;
assign x[2927]= 32'b11110001111000100011111001101100;
assign x[2928]= 32'b11110001111110100011111001110001;
assign x[2929]= 32'b11110010000100110011111001110111;
assign x[2930]= 32'b11110010001010110011111001111100;
assign x[2931]= 32'b11110010010001000011111010000010;
assign x[2932]= 32'b11110010010111000011111010000111;
assign x[2933]= 32'b11110010011101010011111010001100;
assign x[2934]= 32'b11110010100011100011111010010010;
assign x[2935]= 32'b11110010101001100011111010010111;
assign x[2936]= 32'b11110010101111110011111010011100;
assign x[2937]= 32'b11110010110101110011111010100001;
assign x[2938]= 32'b11110010111100000011111010100111;
assign x[2939]= 32'b11110011000010000011111010101100;
assign x[2940]= 32'b11110011001000010011111010110001;
assign x[2941]= 32'b11110011001110100011111010110110;
assign x[2942]= 32'b11110011010100100011111010111011;
assign x[2943]= 32'b11110011011010110011111011000000;
assign x[2944]= 32'b11110011100001000011111011000101;
assign x[2945]= 32'b11110011100111000011111011001010;
assign x[2946]= 32'b11110011101101010011111011001110;
assign x[2947]= 32'b11110011110011100011111011010011;
assign x[2948]= 32'b11110011111001100011111011011000;
assign x[2949]= 32'b11110011111111110011111011011101;
assign x[2950]= 32'b11110100000110000011111011100001;
assign x[2951]= 32'b11110100001100000011111011100110;
assign x[2952]= 32'b11110100010010010011111011101011;
assign x[2953]= 32'b11110100011000100011111011101111;
assign x[2954]= 32'b11110100011110110011111011110100;
assign x[2955]= 32'b11110100100100110011111011111000;
assign x[2956]= 32'b11110100101011000011111011111101;
assign x[2957]= 32'b11110100110001010011111100000001;
assign x[2958]= 32'b11110100110111010011111100000110;
assign x[2959]= 32'b11110100111101100011111100001010;
assign x[2960]= 32'b11110101000011110011111100001110;
assign x[2961]= 32'b11110101001010000011111100010011;
assign x[2962]= 32'b11110101010000000011111100010111;
assign x[2963]= 32'b11110101010110010011111100011011;
assign x[2964]= 32'b11110101011100100011111100011111;
assign x[2965]= 32'b11110101100010110011111100100011;
assign x[2966]= 32'b11110101101001000011111100100111;
assign x[2967]= 32'b11110101101111000011111100101011;
assign x[2968]= 32'b11110101110101010011111100101111;
assign x[2969]= 32'b11110101111011100011111100110011;
assign x[2970]= 32'b11110110000001110011111100110111;
assign x[2971]= 32'b11110110001000000011111100111011;
assign x[2972]= 32'b11110110001110010011111100111111;
assign x[2973]= 32'b11110110010100010011111101000011;
assign x[2974]= 32'b11110110011010100011111101000111;
assign x[2975]= 32'b11110110100000110011111101001010;
assign x[2976]= 32'b11110110100111000011111101001110;
assign x[2977]= 32'b11110110101101010011111101010010;
assign x[2978]= 32'b11110110110011100011111101010101;
assign x[2979]= 32'b11110110111001110011111101011001;
assign x[2980]= 32'b11110110111111110011111101011101;
assign x[2981]= 32'b11110111000110000011111101100000;
assign x[2982]= 32'b11110111001100010011111101100100;
assign x[2983]= 32'b11110111010010100011111101100111;
assign x[2984]= 32'b11110111011000110011111101101010;
assign x[2985]= 32'b11110111011111000011111101101110;
assign x[2986]= 32'b11110111100101010011111101110001;
assign x[2987]= 32'b11110111101011100011111101110100;
assign x[2988]= 32'b11110111110001110011111101111000;
assign x[2989]= 32'b11110111111000000011111101111011;
assign x[2990]= 32'b11110111111110010011111101111110;
assign x[2991]= 32'b11111000000100010011111110000001;
assign x[2992]= 32'b11111000001010100011111110000100;
assign x[2993]= 32'b11111000010000110011111110000111;
assign x[2994]= 32'b11111000010111000011111110001010;
assign x[2995]= 32'b11111000011101010011111110001101;
assign x[2996]= 32'b11111000100011100011111110010000;
assign x[2997]= 32'b11111000101001110011111110010011;
assign x[2998]= 32'b11111000110000000011111110010110;
assign x[2999]= 32'b11111000110110010011111110011001;
assign x[3000]= 32'b11111000111100100011111110011100;
assign x[3001]= 32'b11111001000010110011111110011110;
assign x[3002]= 32'b11111001001001000011111110100001;
assign x[3003]= 32'b11111001001111010011111110100100;
assign x[3004]= 32'b11111001010101100011111110100110;
assign x[3005]= 32'b11111001011011110011111110101001;
assign x[3006]= 32'b11111001100010000011111110101100;
assign x[3007]= 32'b11111001101000010011111110101110;
assign x[3008]= 32'b11111001101110100011111110110001;
assign x[3009]= 32'b11111001110100110011111110110011;
assign x[3010]= 32'b11111001111011000011111110110101;
assign x[3011]= 32'b11111010000001010011111110111000;
assign x[3012]= 32'b11111010000111100011111110111010;
assign x[3013]= 32'b11111010001101110011111110111100;
assign x[3014]= 32'b11111010010100000011111110111111;
assign x[3015]= 32'b11111010011010010011111111000001;
assign x[3016]= 32'b11111010100000100011111111000011;
assign x[3017]= 32'b11111010100110110011111111000101;
assign x[3018]= 32'b11111010101101000011111111000111;
assign x[3019]= 32'b11111010110011010011111111001001;
assign x[3020]= 32'b11111010111001100011111111001011;
assign x[3021]= 32'b11111011000000000011111111001101;
assign x[3022]= 32'b11111011000110010011111111001111;
assign x[3023]= 32'b11111011001100100011111111010001;
assign x[3024]= 32'b11111011010010110011111111010011;
assign x[3025]= 32'b11111011011001000011111111010101;
assign x[3026]= 32'b11111011011111010011111111010111;
assign x[3027]= 32'b11111011100101100011111111011000;
assign x[3028]= 32'b11111011101011110011111111011010;
assign x[3029]= 32'b11111011110010000011111111011100;
assign x[3030]= 32'b11111011111000010011111111011110;
assign x[3031]= 32'b11111011111110100011111111011111;
assign x[3032]= 32'b11111100000100110011111111100001;
assign x[3033]= 32'b11111100001011000011111111100010;
assign x[3034]= 32'b11111100010001010011111111100100;
assign x[3035]= 32'b11111100010111110011111111100101;
assign x[3036]= 32'b11111100011110000011111111100111;
assign x[3037]= 32'b11111100100100010011111111101000;
assign x[3038]= 32'b11111100101010100011111111101001;
assign x[3039]= 32'b11111100110000110011111111101011;
assign x[3040]= 32'b11111100110111000011111111101100;
assign x[3041]= 32'b11111100111101010011111111101101;
assign x[3042]= 32'b11111101000011100011111111101110;
assign x[3043]= 32'b11111101001001110011111111101111;
assign x[3044]= 32'b11111101010000000011111111110000;
assign x[3045]= 32'b11111101010110100011111111110001;
assign x[3046]= 32'b11111101011100110011111111110010;
assign x[3047]= 32'b11111101100011000011111111110011;
assign x[3048]= 32'b11111101101001010011111111110100;
assign x[3049]= 32'b11111101101111100011111111110101;
assign x[3050]= 32'b11111101110101110011111111110110;
assign x[3051]= 32'b11111101111100000011111111110111;
assign x[3052]= 32'b11111110000010010011111111111000;
assign x[3053]= 32'b11111110001000110011111111111001;
assign x[3054]= 32'b11111110001111000011111111111001;
assign x[3055]= 32'b11111110010101010011111111111010;
assign x[3056]= 32'b11111110011011100011111111111011;
assign x[3057]= 32'b11111110100001110011111111111011;
assign x[3058]= 32'b11111110101000000011111111111100;
assign x[3059]= 32'b11111110101110010011111111111100;
assign x[3060]= 32'b11111110110100100011111111111101;
assign x[3061]= 32'b11111110111011000011111111111101;
assign x[3062]= 32'b11111111000001010011111111111110;
assign x[3063]= 32'b11111111000111100011111111111110;
assign x[3064]= 32'b11111111001101110011111111111110;
assign x[3065]= 32'b11111111010100000011111111111111;
assign x[3066]= 32'b11111111011010010011111111111111;
assign x[3067]= 32'b11111111100000100011111111111111;
assign x[3068]= 32'b11111111100110110011111111111111;
assign x[3069]= 32'b11111111101101010011111111111111;
assign x[3070]= 32'b11111111110011100011111111111111;
assign x[3071]= 32'b11111111111001110011111111111111;
assign x[3072]= 32'b11111111111111110100000000000000;
assign x[3073]= 32'b00000000000110010011111111111111;
assign x[3074]= 32'b00000000001100100011111111111111;
assign x[3075]= 32'b00000000010010110011111111111111;
assign x[3076]= 32'b00000000011001000011111111111111;
assign x[3077]= 32'b00000000011111010011111111111111;
assign x[3078]= 32'b00000000100101100011111111111111;
assign x[3079]= 32'b00000000101011110011111111111111;
assign x[3080]= 32'b00000000110010010011111111111110;
assign x[3081]= 32'b00000000111000100011111111111110;
assign x[3082]= 32'b00000000111110110011111111111110;
assign x[3083]= 32'b00000001000101000011111111111101;
assign x[3084]= 32'b00000001001011010011111111111101;
assign x[3085]= 32'b00000001010001100011111111111100;
assign x[3086]= 32'b00000001010111110011111111111100;
assign x[3087]= 32'b00000001011110000011111111111011;
assign x[3088]= 32'b00000001100100100011111111111011;
assign x[3089]= 32'b00000001101010110011111111111010;
assign x[3090]= 32'b00000001110001000011111111111001;
assign x[3091]= 32'b00000001110111010011111111111001;
assign x[3092]= 32'b00000001111101100011111111111000;
assign x[3093]= 32'b00000010000011110011111111110111;
assign x[3094]= 32'b00000010001010000011111111110110;
assign x[3095]= 32'b00000010010000010011111111110101;
assign x[3096]= 32'b00000010010110110011111111110100;
assign x[3097]= 32'b00000010011101000011111111110011;
assign x[3098]= 32'b00000010100011010011111111110010;
assign x[3099]= 32'b00000010101001100011111111110001;
assign x[3100]= 32'b00000010101111110011111111110000;
assign x[3101]= 32'b00000010110110000011111111101111;
assign x[3102]= 32'b00000010111100010011111111101110;
assign x[3103]= 32'b00000011000010100011111111101101;
assign x[3104]= 32'b00000011001000110011111111101100;
assign x[3105]= 32'b00000011001111010011111111101011;
assign x[3106]= 32'b00000011010101100011111111101001;
assign x[3107]= 32'b00000011011011110011111111101000;
assign x[3108]= 32'b00000011100010000011111111100111;
assign x[3109]= 32'b00000011101000010011111111100101;
assign x[3110]= 32'b00000011101110100011111111100100;
assign x[3111]= 32'b00000011110100110011111111100010;
assign x[3112]= 32'b00000011111011000011111111100001;
assign x[3113]= 32'b00000100000001010011111111011111;
assign x[3114]= 32'b00000100000111100011111111011110;
assign x[3115]= 32'b00000100001101110011111111011100;
assign x[3116]= 32'b00000100010100010011111111011010;
assign x[3117]= 32'b00000100011010100011111111011000;
assign x[3118]= 32'b00000100100000110011111111010111;
assign x[3119]= 32'b00000100100111000011111111010101;
assign x[3120]= 32'b00000100101101010011111111010011;
assign x[3121]= 32'b00000100110011100011111111010001;
assign x[3122]= 32'b00000100111001110011111111001111;
assign x[3123]= 32'b00000101000000000011111111001101;
assign x[3124]= 32'b00000101000110010011111111001011;
assign x[3125]= 32'b00000101001100100011111111001001;
assign x[3126]= 32'b00000101010010110011111111000111;
assign x[3127]= 32'b00000101011001000011111111000101;
assign x[3128]= 32'b00000101011111010011111111000011;
assign x[3129]= 32'b00000101100101100011111111000001;
assign x[3130]= 32'b00000101101011110011111110111111;
assign x[3131]= 32'b00000101110010000011111110111100;
assign x[3132]= 32'b00000101111000010011111110111010;
assign x[3133]= 32'b00000101111110100011111110111000;
assign x[3134]= 32'b00000110000100110011111110110101;
assign x[3135]= 32'b00000110001011000011111110110011;
assign x[3136]= 32'b00000110010001010011111110110001;
assign x[3137]= 32'b00000110010111100011111110101110;
assign x[3138]= 32'b00000110011101110011111110101100;
assign x[3139]= 32'b00000110100100000011111110101001;
assign x[3140]= 32'b00000110101010010011111110100110;
assign x[3141]= 32'b00000110110000100011111110100100;
assign x[3142]= 32'b00000110110110110011111110100001;
assign x[3143]= 32'b00000110111101000011111110011110;
assign x[3144]= 32'b00000111000011010011111110011100;
assign x[3145]= 32'b00000111001001100011111110011001;
assign x[3146]= 32'b00000111001111110011111110010110;
assign x[3147]= 32'b00000111010110000011111110010011;
assign x[3148]= 32'b00000111011100010011111110010000;
assign x[3149]= 32'b00000111100010100011111110001101;
assign x[3150]= 32'b00000111101000110011111110001010;
assign x[3151]= 32'b00000111101111000011111110000111;
assign x[3152]= 32'b00000111110101010011111110000100;
assign x[3153]= 32'b00000111111011100011111110000001;
assign x[3154]= 32'b00001000000001110011111101111110;
assign x[3155]= 32'b00001000001000000011111101111011;
assign x[3156]= 32'b00001000001110010011111101111000;
assign x[3157]= 32'b00001000010100100011111101110100;
assign x[3158]= 32'b00001000011010110011111101110001;
assign x[3159]= 32'b00001000100001000011111101101110;
assign x[3160]= 32'b00001000100111000011111101101010;
assign x[3161]= 32'b00001000101101010011111101100111;
assign x[3162]= 32'b00001000110011100011111101100100;
assign x[3163]= 32'b00001000111001110011111101100000;
assign x[3164]= 32'b00001001000000000011111101011101;
assign x[3165]= 32'b00001001000110010011111101011001;
assign x[3166]= 32'b00001001001100100011111101010101;
assign x[3167]= 32'b00001001010010110011111101010010;
assign x[3168]= 32'b00001001011001000011111101001110;
assign x[3169]= 32'b00001001011111000011111101001010;
assign x[3170]= 32'b00001001100101010011111101000111;
assign x[3171]= 32'b00001001101011100011111101000011;
assign x[3172]= 32'b00001001110001110011111100111111;
assign x[3173]= 32'b00001001111000000011111100111011;
assign x[3174]= 32'b00001001111110010011111100110111;
assign x[3175]= 32'b00001010000100010011111100110011;
assign x[3176]= 32'b00001010001010100011111100101111;
assign x[3177]= 32'b00001010010000110011111100101011;
assign x[3178]= 32'b00001010010111000011111100100111;
assign x[3179]= 32'b00001010011101010011111100100011;
assign x[3180]= 32'b00001010100011010011111100011111;
assign x[3181]= 32'b00001010101001100011111100011011;
assign x[3182]= 32'b00001010101111110011111100010111;
assign x[3183]= 32'b00001010110110000011111100010011;
assign x[3184]= 32'b00001010111100010011111100001110;
assign x[3185]= 32'b00001011000010010011111100001010;
assign x[3186]= 32'b00001011001000100011111100000110;
assign x[3187]= 32'b00001011001110110011111100000001;
assign x[3188]= 32'b00001011010101000011111011111101;
assign x[3189]= 32'b00001011011011000011111011111000;
assign x[3190]= 32'b00001011100001010011111011110100;
assign x[3191]= 32'b00001011100111100011111011101111;
assign x[3192]= 32'b00001011101101100011111011101011;
assign x[3193]= 32'b00001011110011110011111011100110;
assign x[3194]= 32'b00001011111010000011111011100001;
assign x[3195]= 32'b00001100000000010011111011011101;
assign x[3196]= 32'b00001100000110010011111011011000;
assign x[3197]= 32'b00001100001100100011111011010011;
assign x[3198]= 32'b00001100010010110011111011001110;
assign x[3199]= 32'b00001100011000110011111011001010;
assign x[3200]= 32'b00001100011111000011111011000101;
assign x[3201]= 32'b00001100100101010011111011000000;
assign x[3202]= 32'b00001100101011010011111010111011;
assign x[3203]= 32'b00001100110001100011111010110110;
assign x[3204]= 32'b00001100110111100011111010110001;
assign x[3205]= 32'b00001100111101110011111010101100;
assign x[3206]= 32'b00001101000100000011111010100111;
assign x[3207]= 32'b00001101001010000011111010100001;
assign x[3208]= 32'b00001101010000010011111010011100;
assign x[3209]= 32'b00001101010110010011111010010111;
assign x[3210]= 32'b00001101011100100011111010010010;
assign x[3211]= 32'b00001101100010110011111010001100;
assign x[3212]= 32'b00001101101000110011111010000111;
assign x[3213]= 32'b00001101101111000011111010000010;
assign x[3214]= 32'b00001101110101000011111001111100;
assign x[3215]= 32'b00001101111011010011111001110111;
assign x[3216]= 32'b00001110000001010011111001110001;
assign x[3217]= 32'b00001110000111100011111001101100;
assign x[3218]= 32'b00001110001101100011111001100110;
assign x[3219]= 32'b00001110010011110011111001100001;
assign x[3220]= 32'b00001110011001110011111001011011;
assign x[3221]= 32'b00001110100000000011111001010101;
assign x[3222]= 32'b00001110100110000011111001010000;
assign x[3223]= 32'b00001110101100010011111001001010;
assign x[3224]= 32'b00001110110010010011111001000100;
assign x[3225]= 32'b00001110111000100011111000111110;
assign x[3226]= 32'b00001110111110100011111000111000;
assign x[3227]= 32'b00001111000100100011111000110011;
assign x[3228]= 32'b00001111001010110011111000101101;
assign x[3229]= 32'b00001111010000110011111000100111;
assign x[3230]= 32'b00001111010111000011111000100001;
assign x[3231]= 32'b00001111011101000011111000011011;
assign x[3232]= 32'b00001111100011000011111000010100;
assign x[3233]= 32'b00001111101001010011111000001110;
assign x[3234]= 32'b00001111101111010011111000001000;
assign x[3235]= 32'b00001111110101100011111000000010;
assign x[3236]= 32'b00001111111011100011110111111100;
assign x[3237]= 32'b00010000000001100011110111110101;
assign x[3238]= 32'b00010000000111110011110111101111;
assign x[3239]= 32'b00010000001101110011110111101001;
assign x[3240]= 32'b00010000010011110011110111100010;
assign x[3241]= 32'b00010000011010000011110111011100;
assign x[3242]= 32'b00010000100000000011110111010110;
assign x[3243]= 32'b00010000100110000011110111001111;
assign x[3244]= 32'b00010000101100000011110111001001;
assign x[3245]= 32'b00010000110010010011110111000010;
assign x[3246]= 32'b00010000111000010011110110111011;
assign x[3247]= 32'b00010000111110010011110110110101;
assign x[3248]= 32'b00010001000100010011110110101110;
assign x[3249]= 32'b00010001001010100011110110100111;
assign x[3250]= 32'b00010001010000100011110110100001;
assign x[3251]= 32'b00010001010110100011110110011010;
assign x[3252]= 32'b00010001011100100011110110010011;
assign x[3253]= 32'b00010001100010100011110110001100;
assign x[3254]= 32'b00010001101000100011110110000101;
assign x[3255]= 32'b00010001101110110011110101111110;
assign x[3256]= 32'b00010001110100110011110101110111;
assign x[3257]= 32'b00010001111010110011110101110000;
assign x[3258]= 32'b00010010000000110011110101101001;
assign x[3259]= 32'b00010010000110110011110101100010;
assign x[3260]= 32'b00010010001100110011110101011011;
assign x[3261]= 32'b00010010010010110011110101010100;
assign x[3262]= 32'b00010010011000110011110101001101;
assign x[3263]= 32'b00010010011110110011110101000101;
assign x[3264]= 32'b00010010100101000011110100111110;
assign x[3265]= 32'b00010010101011000011110100110111;
assign x[3266]= 32'b00010010110001000011110100101111;
assign x[3267]= 32'b00010010110111000011110100101000;
assign x[3268]= 32'b00010010111101000011110100100001;
assign x[3269]= 32'b00010011000011000011110100011001;
assign x[3270]= 32'b00010011001001000011110100010010;
assign x[3271]= 32'b00010011001111000011110100001010;
assign x[3272]= 32'b00010011010101000011110100000010;
assign x[3273]= 32'b00010011011011000011110011111011;
assign x[3274]= 32'b00010011100000110011110011110011;
assign x[3275]= 32'b00010011100110110011110011101100;
assign x[3276]= 32'b00010011101100110011110011100100;
assign x[3277]= 32'b00010011110010110011110011011100;
assign x[3278]= 32'b00010011111000110011110011010100;
assign x[3279]= 32'b00010011111110110011110011001100;
assign x[3280]= 32'b00010100000100110011110011000101;
assign x[3281]= 32'b00010100001010110011110010111101;
assign x[3282]= 32'b00010100010000110011110010110101;
assign x[3283]= 32'b00010100010110100011110010101101;
assign x[3284]= 32'b00010100011100100011110010100101;
assign x[3285]= 32'b00010100100010100011110010011101;
assign x[3286]= 32'b00010100101000100011110010010101;
assign x[3287]= 32'b00010100101110100011110010001100;
assign x[3288]= 32'b00010100110100010011110010000100;
assign x[3289]= 32'b00010100111010010011110001111100;
assign x[3290]= 32'b00010101000000010011110001110100;
assign x[3291]= 32'b00010101000110010011110001101100;
assign x[3292]= 32'b00010101001100000011110001100011;
assign x[3293]= 32'b00010101010010000011110001011011;
assign x[3294]= 32'b00010101011000000011110001010011;
assign x[3295]= 32'b00010101011101110011110001001010;
assign x[3296]= 32'b00010101100011110011110001000010;
assign x[3297]= 32'b00010101101001110011110000111001;
assign x[3298]= 32'b00010101101111100011110000110001;
assign x[3299]= 32'b00010101110101100011110000101000;
assign x[3300]= 32'b00010101111011100011110000100000;
assign x[3301]= 32'b00010110000001010011110000010111;
assign x[3302]= 32'b00010110000111010011110000001110;
assign x[3303]= 32'b00010110001101000011110000000110;
assign x[3304]= 32'b00010110010011000011101111111101;
assign x[3305]= 32'b00010110011001000011101111110100;
assign x[3306]= 32'b00010110011110110011101111101011;
assign x[3307]= 32'b00010110100100110011101111100010;
assign x[3308]= 32'b00010110101010100011101111011010;
assign x[3309]= 32'b00010110110000100011101111010001;
assign x[3310]= 32'b00010110110110010011101111001000;
assign x[3311]= 32'b00010110111100010011101110111111;
assign x[3312]= 32'b00010111000010000011101110110110;
assign x[3313]= 32'b00010111000111110011101110101101;
assign x[3314]= 32'b00010111001101110011101110100011;
assign x[3315]= 32'b00010111010011100011101110011010;
assign x[3316]= 32'b00010111011001100011101110010001;
assign x[3317]= 32'b00010111011111010011101110001000;
assign x[3318]= 32'b00010111100101000011101101111111;
assign x[3319]= 32'b00010111101011000011101101110101;
assign x[3320]= 32'b00010111110000110011101101101100;
assign x[3321]= 32'b00010111110110100011101101100011;
assign x[3322]= 32'b00010111111100100011101101011001;
assign x[3323]= 32'b00011000000010010011101101010000;
assign x[3324]= 32'b00011000001000000011101101000111;
assign x[3325]= 32'b00011000001110000011101100111101;
assign x[3326]= 32'b00011000010011110011101100110100;
assign x[3327]= 32'b00011000011001100011101100101010;
assign x[3328]= 32'b00011000011111010011101100100000;
assign x[3329]= 32'b00011000100101010011101100010111;
assign x[3330]= 32'b00011000101011000011101100001101;
assign x[3331]= 32'b00011000110000110011101100000011;
assign x[3332]= 32'b00011000110110100011101011111010;
assign x[3333]= 32'b00011000111100010011101011110000;
assign x[3334]= 32'b00011001000010000011101011100110;
assign x[3335]= 32'b00011001001000000011101011011100;
assign x[3336]= 32'b00011001001101110011101011010010;
assign x[3337]= 32'b00011001010011100011101011001000;
assign x[3338]= 32'b00011001011001010011101010111110;
assign x[3339]= 32'b00011001011111000011101010110100;
assign x[3340]= 32'b00011001100100110011101010101010;
assign x[3341]= 32'b00011001101010100011101010100000;
assign x[3342]= 32'b00011001110000010011101010010110;
assign x[3343]= 32'b00011001110110000011101010001100;
assign x[3344]= 32'b00011001111011110011101010000010;
assign x[3345]= 32'b00011010000001100011101001111000;
assign x[3346]= 32'b00011010000111010011101001101101;
assign x[3347]= 32'b00011010001101000011101001100011;
assign x[3348]= 32'b00011010010010110011101001011001;
assign x[3349]= 32'b00011010011000100011101001001111;
assign x[3350]= 32'b00011010011110010011101001000100;
assign x[3351]= 32'b00011010100011110011101000111010;
assign x[3352]= 32'b00011010101001100011101000101111;
assign x[3353]= 32'b00011010101111010011101000100101;
assign x[3354]= 32'b00011010110101000011101000011010;
assign x[3355]= 32'b00011010111010110011101000010000;
assign x[3356]= 32'b00011011000000100011101000000101;
assign x[3357]= 32'b00011011000110000011100111111011;
assign x[3358]= 32'b00011011001011110011100111110000;
assign x[3359]= 32'b00011011010001100011100111100101;
assign x[3360]= 32'b00011011010111010011100111011010;
assign x[3361]= 32'b00011011011100110011100111010000;
assign x[3362]= 32'b00011011100010100011100111000101;
assign x[3363]= 32'b00011011101000010011100110111010;
assign x[3364]= 32'b00011011101101110011100110101111;
assign x[3365]= 32'b00011011110011100011100110100100;
assign x[3366]= 32'b00011011111001010011100110011001;
assign x[3367]= 32'b00011011111110110011100110001110;
assign x[3368]= 32'b00011100000100100011100110000011;
assign x[3369]= 32'b00011100001010000011100101111000;
assign x[3370]= 32'b00011100001111110011100101101101;
assign x[3371]= 32'b00011100010101010011100101100010;
assign x[3372]= 32'b00011100011011000011100101010111;
assign x[3373]= 32'b00011100100000110011100101001100;
assign x[3374]= 32'b00011100100110010011100101000001;
assign x[3375]= 32'b00011100101011110011100100110101;
assign x[3376]= 32'b00011100110001100011100100101010;
assign x[3377]= 32'b00011100110111000011100100011111;
assign x[3378]= 32'b00011100111100110011100100010011;
assign x[3379]= 32'b00011101000010010011100100001000;
assign x[3380]= 32'b00011101001000000011100011111101;
assign x[3381]= 32'b00011101001101100011100011110001;
assign x[3382]= 32'b00011101010011000011100011100110;
assign x[3383]= 32'b00011101011000110011100011011010;
assign x[3384]= 32'b00011101011110010011100011001111;
assign x[3385]= 32'b00011101100011110011100011000011;
assign x[3386]= 32'b00011101101001100011100010110111;
assign x[3387]= 32'b00011101101111000011100010101100;
assign x[3388]= 32'b00011101110100100011100010100000;
assign x[3389]= 32'b00011101111010000011100010010100;
assign x[3390]= 32'b00011101111111100011100010001001;
assign x[3391]= 32'b00011110000101010011100001111101;
assign x[3392]= 32'b00011110001010110011100001110001;
assign x[3393]= 32'b00011110010000010011100001100101;
assign x[3394]= 32'b00011110010101110011100001011001;
assign x[3395]= 32'b00011110011011010011100001001101;
assign x[3396]= 32'b00011110100000110011100001000001;
assign x[3397]= 32'b00011110100110010011100000110101;
assign x[3398]= 32'b00011110101100000011100000101001;
assign x[3399]= 32'b00011110110001100011100000011101;
assign x[3400]= 32'b00011110110111000011100000010001;
assign x[3401]= 32'b00011110111100100011100000000101;
assign x[3402]= 32'b00011111000010000011011111111001;
assign x[3403]= 32'b00011111000111100011011111101101;
assign x[3404]= 32'b00011111001101000011011111100000;
assign x[3405]= 32'b00011111010010010011011111010100;
assign x[3406]= 32'b00011111010111110011011111001000;
assign x[3407]= 32'b00011111011101010011011110111011;
assign x[3408]= 32'b00011111100010110011011110101111;
assign x[3409]= 32'b00011111101000010011011110100011;
assign x[3410]= 32'b00011111101101110011011110010110;
assign x[3411]= 32'b00011111110011010011011110001010;
assign x[3412]= 32'b00011111111000100011011101111101;
assign x[3413]= 32'b00011111111110000011011101110001;
assign x[3414]= 32'b00100000000011100011011101100100;
assign x[3415]= 32'b00100000001001000011011101010111;
assign x[3416]= 32'b00100000001110010011011101001011;
assign x[3417]= 32'b00100000010011110011011100111110;
assign x[3418]= 32'b00100000011001010011011100110001;
assign x[3419]= 32'b00100000011110110011011100100101;
assign x[3420]= 32'b00100000100100000011011100011000;
assign x[3421]= 32'b00100000101001100011011100001011;
assign x[3422]= 32'b00100000101110110011011011111110;
assign x[3423]= 32'b00100000110100010011011011110001;
assign x[3424]= 32'b00100000111001110011011011100101;
assign x[3425]= 32'b00100000111111000011011011011000;
assign x[3426]= 32'b00100001000100100011011011001011;
assign x[3427]= 32'b00100001001001110011011010111110;
assign x[3428]= 32'b00100001001111010011011010110001;
assign x[3429]= 32'b00100001010100100011011010100100;
assign x[3430]= 32'b00100001011010000011011010010110;
assign x[3431]= 32'b00100001011111010011011010001001;
assign x[3432]= 32'b00100001100100100011011001111100;
assign x[3433]= 32'b00100001101010000011011001101111;
assign x[3434]= 32'b00100001101111010011011001100010;
assign x[3435]= 32'b00100001110100100011011001010100;
assign x[3436]= 32'b00100001111010000011011001000111;
assign x[3437]= 32'b00100001111111010011011000111010;
assign x[3438]= 32'b00100010000100100011011000101100;
assign x[3439]= 32'b00100010001010000011011000011111;
assign x[3440]= 32'b00100010001111010011011000010010;
assign x[3441]= 32'b00100010010100100011011000000100;
assign x[3442]= 32'b00100010011001110011010111110111;
assign x[3443]= 32'b00100010011111010011010111101001;
assign x[3444]= 32'b00100010100100100011010111011100;
assign x[3445]= 32'b00100010101001110011010111001110;
assign x[3446]= 32'b00100010101111000011010111000000;
assign x[3447]= 32'b00100010110100010011010110110011;
assign x[3448]= 32'b00100010111001100011010110100101;
assign x[3449]= 32'b00100010111110110011010110010111;
assign x[3450]= 32'b00100011000100000011010110001001;
assign x[3451]= 32'b00100011001001010011010101111100;
assign x[3452]= 32'b00100011001110100011010101101110;
assign x[3453]= 32'b00100011010011110011010101100000;
assign x[3454]= 32'b00100011011001000011010101010010;
assign x[3455]= 32'b00100011011110010011010101000100;
assign x[3456]= 32'b00100011100011100011010100110110;
assign x[3457]= 32'b00100011101000110011010100101000;
assign x[3458]= 32'b00100011101110000011010100011010;
assign x[3459]= 32'b00100011110011010011010100001100;
assign x[3460]= 32'b00100011111000010011010011111110;
assign x[3461]= 32'b00100011111101100011010011110000;
assign x[3462]= 32'b00100100000010110011010011100010;
assign x[3463]= 32'b00100100001000000011010011010100;
assign x[3464]= 32'b00100100001101000011010011000110;
assign x[3465]= 32'b00100100010010010011010010110111;
assign x[3466]= 32'b00100100010111100011010010101001;
assign x[3467]= 32'b00100100011100110011010010011011;
assign x[3468]= 32'b00100100100001110011010010001100;
assign x[3469]= 32'b00100100100111000011010001111110;
assign x[3470]= 32'b00100100101100000011010001110000;
assign x[3471]= 32'b00100100110001010011010001100001;
assign x[3472]= 32'b00100100110110100011010001010011;
assign x[3473]= 32'b00100100111011100011010001000100;
assign x[3474]= 32'b00100101000000110011010000110110;
assign x[3475]= 32'b00100101000101110011010000100111;
assign x[3476]= 32'b00100101001011000011010000011001;
assign x[3477]= 32'b00100101010000000011010000001010;
assign x[3478]= 32'b00100101010101000011001111111011;
assign x[3479]= 32'b00100101011010010011001111101101;
assign x[3480]= 32'b00100101011111010011001111011110;
assign x[3481]= 32'b00100101100100100011001111001111;
assign x[3482]= 32'b00100101101001100011001111000001;
assign x[3483]= 32'b00100101101110100011001110110010;
assign x[3484]= 32'b00100101110011110011001110100011;
assign x[3485]= 32'b00100101111000110011001110010100;
assign x[3486]= 32'b00100101111101110011001110000101;
assign x[3487]= 32'b00100110000010110011001101110110;
assign x[3488]= 32'b00100110000111110011001101100111;
assign x[3489]= 32'b00100110001101000011001101011000;
assign x[3490]= 32'b00100110010010000011001101001001;
assign x[3491]= 32'b00100110010111000011001100111010;
assign x[3492]= 32'b00100110011100000011001100101011;
assign x[3493]= 32'b00100110100001000011001100011100;
assign x[3494]= 32'b00100110100110000011001100001101;
assign x[3495]= 32'b00100110101011000011001011111110;
assign x[3496]= 32'b00100110110000000011001011101110;
assign x[3497]= 32'b00100110110101000011001011011111;
assign x[3498]= 32'b00100110111010000011001011010000;
assign x[3499]= 32'b00100110111111000011001011000001;
assign x[3500]= 32'b00100111000100000011001010110001;
assign x[3501]= 32'b00100111001001000011001010100010;
assign x[3502]= 32'b00100111001110000011001010010011;
assign x[3503]= 32'b00100111010011000011001010000011;
assign x[3504]= 32'b00100111010111110011001001110100;
assign x[3505]= 32'b00100111011100110011001001100100;
assign x[3506]= 32'b00100111100001110011001001010101;
assign x[3507]= 32'b00100111100110110011001001000101;
assign x[3508]= 32'b00100111101011110011001000110110;
assign x[3509]= 32'b00100111110000100011001000100110;
assign x[3510]= 32'b00100111110101100011001000010110;
assign x[3511]= 32'b00100111111010100011001000000111;
assign x[3512]= 32'b00100111111111010011000111110111;
assign x[3513]= 32'b00101000000100010011000111100111;
assign x[3514]= 32'b00101000001001000011000111011000;
assign x[3515]= 32'b00101000001110000011000111001000;
assign x[3516]= 32'b00101000010010110011000110111000;
assign x[3517]= 32'b00101000010111110011000110101000;
assign x[3518]= 32'b00101000011100100011000110011000;
assign x[3519]= 32'b00101000100001100011000110001000;
assign x[3520]= 32'b00101000100110010011000101111001;
assign x[3521]= 32'b00101000101011010011000101101001;
assign x[3522]= 32'b00101000110000000011000101011001;
assign x[3523]= 32'b00101000110101000011000101001001;
assign x[3524]= 32'b00101000111001110011000100111000;
assign x[3525]= 32'b00101000111110100011000100101000;
assign x[3526]= 32'b00101001000011100011000100011000;
assign x[3527]= 32'b00101001001000010011000100001000;
assign x[3528]= 32'b00101001001101000011000011111000;
assign x[3529]= 32'b00101001010001110011000011101000;
assign x[3530]= 32'b00101001010110100011000011011000;
assign x[3531]= 32'b00101001011011100011000011000111;
assign x[3532]= 32'b00101001100000010011000010110111;
assign x[3533]= 32'b00101001100101000011000010100111;
assign x[3534]= 32'b00101001101001110011000010010110;
assign x[3535]= 32'b00101001101110100011000010000110;
assign x[3536]= 32'b00101001110011010011000001110110;
assign x[3537]= 32'b00101001111000000011000001100101;
assign x[3538]= 32'b00101001111100110011000001010101;
assign x[3539]= 32'b00101010000001100011000001000100;
assign x[3540]= 32'b00101010000110010011000000110100;
assign x[3541]= 32'b00101010001011000011000000100011;
assign x[3542]= 32'b00101010001111110011000000010011;
assign x[3543]= 32'b00101010010100100011000000000010;
assign x[3544]= 32'b00101010011001010010111111110001;
assign x[3545]= 32'b00101010011101110010111111100001;
assign x[3546]= 32'b00101010100010100010111111010000;
assign x[3547]= 32'b00101010100111010010111110111111;
assign x[3548]= 32'b00101010101100000010111110101111;
assign x[3549]= 32'b00101010110000100010111110011110;
assign x[3550]= 32'b00101010110101010010111110001101;
assign x[3551]= 32'b00101010111010000010111101111100;
assign x[3552]= 32'b00101010111110100010111101101011;
assign x[3553]= 32'b00101011000011010010111101011010;
assign x[3554]= 32'b00101011001000000010111101001001;
assign x[3555]= 32'b00101011001100100010111100111000;
assign x[3556]= 32'b00101011010001010010111100101000;
assign x[3557]= 32'b00101011010101110010111100010110;
assign x[3558]= 32'b00101011011010100010111100000101;
assign x[3559]= 32'b00101011011111000010111011110100;
assign x[3560]= 32'b00101011100011100010111011100011;
assign x[3561]= 32'b00101011101000010010111011010010;
assign x[3562]= 32'b00101011101100110010111011000001;
assign x[3563]= 32'b00101011110001100010111010110000;
assign x[3564]= 32'b00101011110110000010111010011111;
assign x[3565]= 32'b00101011111010100010111010001101;
assign x[3566]= 32'b00101011111111000010111001111100;
assign x[3567]= 32'b00101100000011110010111001101011;
assign x[3568]= 32'b00101100001000010010111001011010;
assign x[3569]= 32'b00101100001100110010111001001000;
assign x[3570]= 32'b00101100010001010010111000110111;
assign x[3571]= 32'b00101100010101110010111000100101;
assign x[3572]= 32'b00101100011010100010111000010100;
assign x[3573]= 32'b00101100011111000010111000000011;
assign x[3574]= 32'b00101100100011100010110111110001;
assign x[3575]= 32'b00101100101000000010110111100000;
assign x[3576]= 32'b00101100101100100010110111001110;
assign x[3577]= 32'b00101100110001000010110110111100;
assign x[3578]= 32'b00101100110101100010110110101011;
assign x[3579]= 32'b00101100111010000010110110011001;
assign x[3580]= 32'b00101100111110010010110110001000;
assign x[3581]= 32'b00101101000010110010110101110110;
assign x[3582]= 32'b00101101000111010010110101100100;
assign x[3583]= 32'b00101101001011110010110101010010;
assign x[3584]= 32'b00101101010000010010110101000001;
assign x[3585]= 32'b00101101010100100010110100101111;
assign x[3586]= 32'b00101101011001000010110100011101;
assign x[3587]= 32'b00101101011101100010110100001011;
assign x[3588]= 32'b00101101100010000010110011111001;
assign x[3589]= 32'b00101101100110010010110011101000;
assign x[3590]= 32'b00101101101010110010110011010110;
assign x[3591]= 32'b00101101101111000010110011000100;
assign x[3592]= 32'b00101101110011100010110010110010;
assign x[3593]= 32'b00101101111000000010110010100000;
assign x[3594]= 32'b00101101111100010010110010001110;
assign x[3595]= 32'b00101110000000110010110001111100;
assign x[3596]= 32'b00101110000101000010110001101010;
assign x[3597]= 32'b00101110001001010010110001010111;
assign x[3598]= 32'b00101110001101110010110001000101;
assign x[3599]= 32'b00101110010010000010110000110011;
assign x[3600]= 32'b00101110010110100010110000100001;
assign x[3601]= 32'b00101110011010110010110000001111;
assign x[3602]= 32'b00101110011111000010101111111100;
assign x[3603]= 32'b00101110100011010010101111101010;
assign x[3604]= 32'b00101110100111110010101111011000;
assign x[3605]= 32'b00101110101100000010101111000110;
assign x[3606]= 32'b00101110110000010010101110110011;
assign x[3607]= 32'b00101110110100100010101110100001;
assign x[3608]= 32'b00101110111000110010101110001110;
assign x[3609]= 32'b00101110111101000010101101111100;
assign x[3610]= 32'b00101111000001010010101101101010;
assign x[3611]= 32'b00101111000101100010101101010111;
assign x[3612]= 32'b00101111001010000010101101000101;
assign x[3613]= 32'b00101111001110000010101100110010;
assign x[3614]= 32'b00101111010010010010101100100000;
assign x[3615]= 32'b00101111010110100010101100001101;
assign x[3616]= 32'b00101111011010110010101011111010;
assign x[3617]= 32'b00101111011111000010101011101000;
assign x[3618]= 32'b00101111100011010010101011010101;
assign x[3619]= 32'b00101111100111100010101011000010;
assign x[3620]= 32'b00101111101011110010101010110000;
assign x[3621]= 32'b00101111101111110010101010011101;
assign x[3622]= 32'b00101111110100000010101010001010;
assign x[3623]= 32'b00101111111000010010101001110111;
assign x[3624]= 32'b00101111111100010010101001100101;
assign x[3625]= 32'b00110000000000100010101001010010;
assign x[3626]= 32'b00110000000100110010101000111111;
assign x[3627]= 32'b00110000001000110010101000101100;
assign x[3628]= 32'b00110000001101000010101000011001;
assign x[3629]= 32'b00110000010001000010101000000110;
assign x[3630]= 32'b00110000010101010010100111110011;
assign x[3631]= 32'b00110000011001010010100111100000;
assign x[3632]= 32'b00110000011101100010100111001101;
assign x[3633]= 32'b00110000100001100010100110111010;
assign x[3634]= 32'b00110000100101100010100110100111;
assign x[3635]= 32'b00110000101001110010100110010100;
assign x[3636]= 32'b00110000101101110010100110000001;
assign x[3637]= 32'b00110000110001110010100101101110;
assign x[3638]= 32'b00110000110110000010100101011010;
assign x[3639]= 32'b00110000111010000010100101000111;
assign x[3640]= 32'b00110000111110000010100100110100;
assign x[3641]= 32'b00110001000010000010100100100001;
assign x[3642]= 32'b00110001000110000010100100001110;
assign x[3643]= 32'b00110001001010000010100011111010;
assign x[3644]= 32'b00110001001110000010100011100111;
assign x[3645]= 32'b00110001010010010010100011010100;
assign x[3646]= 32'b00110001010110010010100011000000;
assign x[3647]= 32'b00110001011010010010100010101101;
assign x[3648]= 32'b00110001011110010010100010011001;
assign x[3649]= 32'b00110001100010000010100010000110;
assign x[3650]= 32'b00110001100110000010100001110010;
assign x[3651]= 32'b00110001101010000010100001011111;
assign x[3652]= 32'b00110001101110000010100001001011;
assign x[3653]= 32'b00110001110010000010100000111000;
assign x[3654]= 32'b00110001110110000010100000100100;
assign x[3655]= 32'b00110001111001110010100000010001;
assign x[3656]= 32'b00110001111101110010011111111101;
assign x[3657]= 32'b00110010000001110010011111101010;
assign x[3658]= 32'b00110010000101100010011111010110;
assign x[3659]= 32'b00110010001001100010011111000010;
assign x[3660]= 32'b00110010001101100010011110101111;
assign x[3661]= 32'b00110010010001010010011110011011;
assign x[3662]= 32'b00110010010101010010011110000111;
assign x[3663]= 32'b00110010011001000010011101110011;
assign x[3664]= 32'b00110010011101000010011101011111;
assign x[3665]= 32'b00110010100000110010011101001100;
assign x[3666]= 32'b00110010100100110010011100111000;
assign x[3667]= 32'b00110010101000100010011100100100;
assign x[3668]= 32'b00110010101100010010011100010000;
assign x[3669]= 32'b00110010110000010010011011111100;
assign x[3670]= 32'b00110010110100000010011011101000;
assign x[3671]= 32'b00110010110111110010011011010100;
assign x[3672]= 32'b00110010111011100010011011000000;
assign x[3673]= 32'b00110010111111100010011010101100;
assign x[3674]= 32'b00110011000011010010011010011000;
assign x[3675]= 32'b00110011000111000010011010000100;
assign x[3676]= 32'b00110011001010110010011001110000;
assign x[3677]= 32'b00110011001110100010011001011100;
assign x[3678]= 32'b00110011010010010010011001001000;
assign x[3679]= 32'b00110011010110000010011000110100;
assign x[3680]= 32'b00110011011001110010011000011111;
assign x[3681]= 32'b00110011011101100010011000001011;
assign x[3682]= 32'b00110011100001010010010111110111;
assign x[3683]= 32'b00110011100101000010010111100011;
assign x[3684]= 32'b00110011101000110010010111001111;
assign x[3685]= 32'b00110011101100100010010110111010;
assign x[3686]= 32'b00110011110000010010010110100110;
assign x[3687]= 32'b00110011110011110010010110010010;
assign x[3688]= 32'b00110011110111100010010101111101;
assign x[3689]= 32'b00110011111011010010010101101001;
assign x[3690]= 32'b00110011111110110010010101010100;
assign x[3691]= 32'b00110100000010100010010101000000;
assign x[3692]= 32'b00110100000110010010010100101100;
assign x[3693]= 32'b00110100001001110010010100010111;
assign x[3694]= 32'b00110100001101100010010100000011;
assign x[3695]= 32'b00110100010001000010010011101110;
assign x[3696]= 32'b00110100010100110010010011011010;
assign x[3697]= 32'b00110100011000010010010011000101;
assign x[3698]= 32'b00110100011100000010010010110000;
assign x[3699]= 32'b00110100011111100010010010011100;
assign x[3700]= 32'b00110100100011000010010010000111;
assign x[3701]= 32'b00110100100110110010010001110011;
assign x[3702]= 32'b00110100101010010010010001011110;
assign x[3703]= 32'b00110100101101110010010001001001;
assign x[3704]= 32'b00110100110001100010010000110100;
assign x[3705]= 32'b00110100110101000010010000100000;
assign x[3706]= 32'b00110100111000100010010000001011;
assign x[3707]= 32'b00110100111100000010001111110110;
assign x[3708]= 32'b00110100111111100010001111100001;
assign x[3709]= 32'b00110101000011000010001111001101;
assign x[3710]= 32'b00110101000110100010001110111000;
assign x[3711]= 32'b00110101001010000010001110100011;
assign x[3712]= 32'b00110101001101100010001110001110;
assign x[3713]= 32'b00110101010001000010001101111001;
assign x[3714]= 32'b00110101010100100010001101100100;
assign x[3715]= 32'b00110101011000000010001101001111;
assign x[3716]= 32'b00110101011011100010001100111010;
assign x[3717]= 32'b00110101011111000010001100100101;
assign x[3718]= 32'b00110101100010010010001100010000;
assign x[3719]= 32'b00110101100101110010001011111011;
assign x[3720]= 32'b00110101101001010010001011100110;
assign x[3721]= 32'b00110101101100110010001011010001;
assign x[3722]= 32'b00110101110000000010001010111100;
assign x[3723]= 32'b00110101110011100010001010100111;
assign x[3724]= 32'b00110101110111000010001010010010;
assign x[3725]= 32'b00110101111010010010001001111101;
assign x[3726]= 32'b00110101111101110010001001100111;
assign x[3727]= 32'b00110110000001000010001001010010;
assign x[3728]= 32'b00110110000100100010001000111101;
assign x[3729]= 32'b00110110000111110010001000101000;
assign x[3730]= 32'b00110110001011000010001000010010;
assign x[3731]= 32'b00110110001110100010000111111101;
assign x[3732]= 32'b00110110010001110010000111101000;
assign x[3733]= 32'b00110110010101000010000111010010;
assign x[3734]= 32'b00110110011000100010000110111101;
assign x[3735]= 32'b00110110011011110010000110101000;
assign x[3736]= 32'b00110110011111000010000110010010;
assign x[3737]= 32'b00110110100010010010000101111101;
assign x[3738]= 32'b00110110100101100010000101101000;
assign x[3739]= 32'b00110110101001000010000101010010;
assign x[3740]= 32'b00110110101100010010000100111101;
assign x[3741]= 32'b00110110101111100010000100100111;
assign x[3742]= 32'b00110110110010110010000100010010;
assign x[3743]= 32'b00110110110110000010000011111100;
assign x[3744]= 32'b00110110111001010010000011100111;
assign x[3745]= 32'b00110110111100010010000011010001;
assign x[3746]= 32'b00110110111111100010000010111011;
assign x[3747]= 32'b00110111000010110010000010100110;
assign x[3748]= 32'b00110111000110000010000010010000;
assign x[3749]= 32'b00110111001001010010000001111011;
assign x[3750]= 32'b00110111001100010010000001100101;
assign x[3751]= 32'b00110111001111100010000001001111;
assign x[3752]= 32'b00110111010010110010000000111001;
assign x[3753]= 32'b00110111010101110010000000100100;
assign x[3754]= 32'b00110111011001000010000000001110;
assign x[3755]= 32'b00110111011100010001111111111000;
assign x[3756]= 32'b00110111011111010001111111100010;
assign x[3757]= 32'b00110111100010100001111111001101;
assign x[3758]= 32'b00110111100101100001111110110111;
assign x[3759]= 32'b00110111101000110001111110100001;
assign x[3760]= 32'b00110111101011110001111110001011;
assign x[3761]= 32'b00110111101110110001111101110101;
assign x[3762]= 32'b00110111110010000001111101011111;
assign x[3763]= 32'b00110111110101000001111101001001;
assign x[3764]= 32'b00110111111000000001111100110100;
assign x[3765]= 32'b00110111111011010001111100011110;
assign x[3766]= 32'b00110111111110010001111100001000;
assign x[3767]= 32'b00111000000001010001111011110010;
assign x[3768]= 32'b00111000000100010001111011011100;
assign x[3769]= 32'b00111000000111010001111011000110;
assign x[3770]= 32'b00111000001010010001111010110000;
assign x[3771]= 32'b00111000001101010001111010011001;
assign x[3772]= 32'b00111000010000010001111010000011;
assign x[3773]= 32'b00111000010011010001111001101101;
assign x[3774]= 32'b00111000010110010001111001010111;
assign x[3775]= 32'b00111000011001010001111001000001;
assign x[3776]= 32'b00111000011100010001111000101011;
assign x[3777]= 32'b00111000011111010001111000010101;
assign x[3778]= 32'b00111000100010010001110111111110;
assign x[3779]= 32'b00111000100101000001110111101000;
assign x[3780]= 32'b00111000101000000001110111010010;
assign x[3781]= 32'b00111000101011000001110110111100;
assign x[3782]= 32'b00111000101101110001110110100110;
assign x[3783]= 32'b00111000110000110001110110001111;
assign x[3784]= 32'b00111000110011110001110101111001;
assign x[3785]= 32'b00111000110110100001110101100011;
assign x[3786]= 32'b00111000111001100001110101001100;
assign x[3787]= 32'b00111000111100010001110100110110;
assign x[3788]= 32'b00111000111111010001110100100000;
assign x[3789]= 32'b00111001000010000001110100001001;
assign x[3790]= 32'b00111001000100110001110011110011;
assign x[3791]= 32'b00111001000111110001110011011100;
assign x[3792]= 32'b00111001001010100001110011000110;
assign x[3793]= 32'b00111001001101010001110010101111;
assign x[3794]= 32'b00111001010000010001110010011001;
assign x[3795]= 32'b00111001010011000001110010000011;
assign x[3796]= 32'b00111001010101110001110001101100;
assign x[3797]= 32'b00111001011000100001110001010101;
assign x[3798]= 32'b00111001011011010001110000111111;
assign x[3799]= 32'b00111001011110000001110000101000;
assign x[3800]= 32'b00111001100000110001110000010010;
assign x[3801]= 32'b00111001100011100001101111111011;
assign x[3802]= 32'b00111001100110010001101111100101;
assign x[3803]= 32'b00111001101001000001101111001110;
assign x[3804]= 32'b00111001101011110001101110110111;
assign x[3805]= 32'b00111001101110100001101110100001;
assign x[3806]= 32'b00111001110001010001101110001010;
assign x[3807]= 32'b00111001110100000001101101110011;
assign x[3808]= 32'b00111001110110100001101101011101;
assign x[3809]= 32'b00111001111001010001101101000110;
assign x[3810]= 32'b00111001111100000001101100101111;
assign x[3811]= 32'b00111001111110110001101100011000;
assign x[3812]= 32'b00111010000001010001101100000010;
assign x[3813]= 32'b00111010000100000001101011101011;
assign x[3814]= 32'b00111010000110100001101011010100;
assign x[3815]= 32'b00111010001001010001101010111101;
assign x[3816]= 32'b00111010001011110001101010100110;
assign x[3817]= 32'b00111010001110100001101010001111;
assign x[3818]= 32'b00111010010001000001101001111001;
assign x[3819]= 32'b00111010010011110001101001100010;
assign x[3820]= 32'b00111010010110010001101001001011;
assign x[3821]= 32'b00111010011000110001101000110100;
assign x[3822]= 32'b00111010011011010001101000011101;
assign x[3823]= 32'b00111010011110000001101000000110;
assign x[3824]= 32'b00111010100000100001100111101111;
assign x[3825]= 32'b00111010100011000001100111011000;
assign x[3826]= 32'b00111010100101100001100111000001;
assign x[3827]= 32'b00111010101000000001100110101010;
assign x[3828]= 32'b00111010101010100001100110010011;
assign x[3829]= 32'b00111010101101000001100101111100;
assign x[3830]= 32'b00111010101111100001100101100101;
assign x[3831]= 32'b00111010110010000001100101001110;
assign x[3832]= 32'b00111010110100100001100100110111;
assign x[3833]= 32'b00111010110111000001100100100000;
assign x[3834]= 32'b00111010111001100001100100001000;
assign x[3835]= 32'b00111010111100000001100011110001;
assign x[3836]= 32'b00111010111110100001100011011010;
assign x[3837]= 32'b00111011000000110001100011000011;
assign x[3838]= 32'b00111011000011010001100010101100;
assign x[3839]= 32'b00111011000101110001100010010101;
assign x[3840]= 32'b00111011001000000001100001111101;
assign x[3841]= 32'b00111011001010100001100001100110;
assign x[3842]= 32'b00111011001101000001100001001111;
assign x[3843]= 32'b00111011001111010001100000111000;
assign x[3844]= 32'b00111011010001110001100000100000;
assign x[3845]= 32'b00111011010100000001100000001001;
assign x[3846]= 32'b00111011010110010001011111110010;
assign x[3847]= 32'b00111011011000110001011111011010;
assign x[3848]= 32'b00111011011011000001011111000011;
assign x[3849]= 32'b00111011011101010001011110101100;
assign x[3850]= 32'b00111011011111110001011110010100;
assign x[3851]= 32'b00111011100010000001011101111101;
assign x[3852]= 32'b00111011100100010001011101100110;
assign x[3853]= 32'b00111011100110100001011101001110;
assign x[3854]= 32'b00111011101000110001011100110111;
assign x[3855]= 32'b00111011101011010001011100011111;
assign x[3856]= 32'b00111011101101100001011100001000;
assign x[3857]= 32'b00111011101111110001011011110001;
assign x[3858]= 32'b00111011110010000001011011011001;
assign x[3859]= 32'b00111011110100010001011011000010;
assign x[3860]= 32'b00111011110110100001011010101010;
assign x[3861]= 32'b00111011111000100001011010010011;
assign x[3862]= 32'b00111011111010110001011001111011;
assign x[3863]= 32'b00111011111101000001011001100100;
assign x[3864]= 32'b00111011111111010001011001001100;
assign x[3865]= 32'b00111100000001100001011000110100;
assign x[3866]= 32'b00111100000011100001011000011101;
assign x[3867]= 32'b00111100000101110001011000000101;
assign x[3868]= 32'b00111100001000000001010111101110;
assign x[3869]= 32'b00111100001010000001010111010110;
assign x[3870]= 32'b00111100001100010001010110111110;
assign x[3871]= 32'b00111100001110010001010110100111;
assign x[3872]= 32'b00111100010000100001010110001111;
assign x[3873]= 32'b00111100010010100001010101110111;
assign x[3874]= 32'b00111100010100110001010101100000;
assign x[3875]= 32'b00111100010110110001010101001000;
assign x[3876]= 32'b00111100011000110001010100110000;
assign x[3877]= 32'b00111100011011000001010100011001;
assign x[3878]= 32'b00111100011101000001010100000001;
assign x[3879]= 32'b00111100011111000001010011101001;
assign x[3880]= 32'b00111100100001000001010011010001;
assign x[3881]= 32'b00111100100011000001010010111010;
assign x[3882]= 32'b00111100100101010001010010100010;
assign x[3883]= 32'b00111100100111010001010010001010;
assign x[3884]= 32'b00111100101001010001010001110010;
assign x[3885]= 32'b00111100101011010001010001011010;
assign x[3886]= 32'b00111100101101010001010001000011;
assign x[3887]= 32'b00111100101111010001010000101011;
assign x[3888]= 32'b00111100110001010001010000010011;
assign x[3889]= 32'b00111100110011000001001111111011;
assign x[3890]= 32'b00111100110101000001001111100011;
assign x[3891]= 32'b00111100110111000001001111001011;
assign x[3892]= 32'b00111100111001000001001110110011;
assign x[3893]= 32'b00111100111011000001001110011011;
assign x[3894]= 32'b00111100111100110001001110000011;
assign x[3895]= 32'b00111100111110110001001101101100;
assign x[3896]= 32'b00111101000000100001001101010100;
assign x[3897]= 32'b00111101000010100001001100111100;
assign x[3898]= 32'b00111101000100100001001100100100;
assign x[3899]= 32'b00111101000110010001001100001100;
assign x[3900]= 32'b00111101001000010001001011110100;
assign x[3901]= 32'b00111101001010000001001011011100;
assign x[3902]= 32'b00111101001011110001001011000100;
assign x[3903]= 32'b00111101001101110001001010101100;
assign x[3904]= 32'b00111101001111100001001010010100;
assign x[3905]= 32'b00111101010001010001001001111011;
assign x[3906]= 32'b00111101010011010001001001100011;
assign x[3907]= 32'b00111101010101000001001001001011;
assign x[3908]= 32'b00111101010110110001001000110011;
assign x[3909]= 32'b00111101011000100001001000011011;
assign x[3910]= 32'b00111101011010010001001000000011;
assign x[3911]= 32'b00111101011100000001000111101011;
assign x[3912]= 32'b00111101011101110001000111010011;
assign x[3913]= 32'b00111101011111100001000110111011;
assign x[3914]= 32'b00111101100001010001000110100010;
assign x[3915]= 32'b00111101100011000001000110001010;
assign x[3916]= 32'b00111101100100110001000101110010;
assign x[3917]= 32'b00111101100110100001000101011010;
assign x[3918]= 32'b00111101101000010001000101000010;
assign x[3919]= 32'b00111101101001110001000100101010;
assign x[3920]= 32'b00111101101011100001000100010001;
assign x[3921]= 32'b00111101101101010001000011111001;
assign x[3922]= 32'b00111101101110110001000011100001;
assign x[3923]= 32'b00111101110000100001000011001001;
assign x[3924]= 32'b00111101110010010001000010110000;
assign x[3925]= 32'b00111101110011110001000010011000;
assign x[3926]= 32'b00111101110101100001000010000000;
assign x[3927]= 32'b00111101110111000001000001101000;
assign x[3928]= 32'b00111101111000100001000001001111;
assign x[3929]= 32'b00111101111010010001000000110111;
assign x[3930]= 32'b00111101111011110001000000011111;
assign x[3931]= 32'b00111101111101010001000000000110;
assign x[3932]= 32'b00111101111111000000111111101110;
assign x[3933]= 32'b00111110000000100000111111010110;
assign x[3934]= 32'b00111110000010000000111110111101;
assign x[3935]= 32'b00111110000011100000111110100101;
assign x[3936]= 32'b00111110000101000000111110001100;
assign x[3937]= 32'b00111110000110110000111101110100;
assign x[3938]= 32'b00111110001000010000111101011100;
assign x[3939]= 32'b00111110001001110000111101000011;
assign x[3940]= 32'b00111110001011010000111100101011;
assign x[3941]= 32'b00111110001100110000111100010010;
assign x[3942]= 32'b00111110001110000000111011111010;
assign x[3943]= 32'b00111110001111100000111011100010;
assign x[3944]= 32'b00111110010001000000111011001001;
assign x[3945]= 32'b00111110010010100000111010110001;
assign x[3946]= 32'b00111110010100000000111010011000;
assign x[3947]= 32'b00111110010101010000111010000000;
assign x[3948]= 32'b00111110010110110000111001100111;
assign x[3949]= 32'b00111110011000010000111001001111;
assign x[3950]= 32'b00111110011001100000111000110110;
assign x[3951]= 32'b00111110011011000000111000011110;
assign x[3952]= 32'b00111110011100010000111000000101;
assign x[3953]= 32'b00111110011101110000110111101101;
assign x[3954]= 32'b00111110011111000000110111010100;
assign x[3955]= 32'b00111110100000100000110110111100;
assign x[3956]= 32'b00111110100001110000110110100011;
assign x[3957]= 32'b00111110100011000000110110001011;
assign x[3958]= 32'b00111110100100100000110101110010;
assign x[3959]= 32'b00111110100101110000110101011001;
assign x[3960]= 32'b00111110100111000000110101000001;
assign x[3961]= 32'b00111110101000010000110100101000;
assign x[3962]= 32'b00111110101001110000110100010000;
assign x[3963]= 32'b00111110101011000000110011110111;
assign x[3964]= 32'b00111110101100010000110011011110;
assign x[3965]= 32'b00111110101101100000110011000110;
assign x[3966]= 32'b00111110101110110000110010101101;
assign x[3967]= 32'b00111110110000000000110010010101;
assign x[3968]= 32'b00111110110001010000110001111100;
assign x[3969]= 32'b00111110110010100000110001100011;
assign x[3970]= 32'b00111110110011100000110001001011;
assign x[3971]= 32'b00111110110100110000110000110010;
assign x[3972]= 32'b00111110110110000000110000011001;
assign x[3973]= 32'b00111110110111010000110000000001;
assign x[3974]= 32'b00111110111000010000101111101000;
assign x[3975]= 32'b00111110111001100000101111001111;
assign x[3976]= 32'b00111110111010110000101110110110;
assign x[3977]= 32'b00111110111011110000101110011110;
assign x[3978]= 32'b00111110111101000000101110000101;
assign x[3979]= 32'b00111110111110000000101101101100;
assign x[3980]= 32'b00111110111111010000101101010100;
assign x[3981]= 32'b00111111000000010000101100111011;
assign x[3982]= 32'b00111111000001100000101100100010;
assign x[3983]= 32'b00111111000010100000101100001001;
assign x[3984]= 32'b00111111000011100000101011110001;
assign x[3985]= 32'b00111111000100110000101011011000;
assign x[3986]= 32'b00111111000101110000101010111111;
assign x[3987]= 32'b00111111000110110000101010100110;
assign x[3988]= 32'b00111111000111110000101010001101;
assign x[3989]= 32'b00111111001000110000101001110101;
assign x[3990]= 32'b00111111001001110000101001011100;
assign x[3991]= 32'b00111111001010110000101001000011;
assign x[3992]= 32'b00111111001011110000101000101010;
assign x[3993]= 32'b00111111001100110000101000010001;
assign x[3994]= 32'b00111111001101110000100111111001;
assign x[3995]= 32'b00111111001110110000100111100000;
assign x[3996]= 32'b00111111001111110000100111000111;
assign x[3997]= 32'b00111111010000110000100110101110;
assign x[3998]= 32'b00111111010001110000100110010101;
assign x[3999]= 32'b00111111010010100000100101111100;
assign x[4000]= 32'b00111111010011100000100101100100;
assign x[4001]= 32'b00111111010100100000100101001011;
assign x[4002]= 32'b00111111010101010000100100110010;
assign x[4003]= 32'b00111111010110010000100100011001;
assign x[4004]= 32'b00111111010111010000100100000000;
assign x[4005]= 32'b00111111011000000000100011100111;
assign x[4006]= 32'b00111111011001000000100011001110;
assign x[4007]= 32'b00111111011001110000100010110101;
assign x[4008]= 32'b00111111011010100000100010011100;
assign x[4009]= 32'b00111111011011100000100010000100;
assign x[4010]= 32'b00111111011100010000100001101011;
assign x[4011]= 32'b00111111011101000000100001010010;
assign x[4012]= 32'b00111111011110000000100000111001;
assign x[4013]= 32'b00111111011110110000100000100000;
assign x[4014]= 32'b00111111011111100000100000000111;
assign x[4015]= 32'b00111111100000010000011111101110;
assign x[4016]= 32'b00111111100001000000011111010101;
assign x[4017]= 32'b00111111100001110000011110111100;
assign x[4018]= 32'b00111111100010100000011110100011;
assign x[4019]= 32'b00111111100011010000011110001010;
assign x[4020]= 32'b00111111100100000000011101110001;
assign x[4021]= 32'b00111111100100110000011101011000;
assign x[4022]= 32'b00111111100101100000011100111111;
assign x[4023]= 32'b00111111100110010000011100100110;
assign x[4024]= 32'b00111111100111000000011100001101;
assign x[4025]= 32'b00111111100111100000011011110100;
assign x[4026]= 32'b00111111101000010000011011011011;
assign x[4027]= 32'b00111111101001000000011011000010;
assign x[4028]= 32'b00111111101001100000011010101001;
assign x[4029]= 32'b00111111101010010000011010010000;
assign x[4030]= 32'b00111111101011000000011001110111;
assign x[4031]= 32'b00111111101011100000011001011110;
assign x[4032]= 32'b00111111101100010000011001000101;
assign x[4033]= 32'b00111111101100110000011000101100;
assign x[4034]= 32'b00111111101101010000011000010011;
assign x[4035]= 32'b00111111101110000000010111111010;
assign x[4036]= 32'b00111111101110100000010111100001;
assign x[4037]= 32'b00111111101111000000010111001000;
assign x[4038]= 32'b00111111101111110000010110101111;
assign x[4039]= 32'b00111111110000010000010110010110;
assign x[4040]= 32'b00111111110000110000010101111101;
assign x[4041]= 32'b00111111110001010000010101100100;
assign x[4042]= 32'b00111111110001110000010101001011;
assign x[4043]= 32'b00111111110010010000010100110010;
assign x[4044]= 32'b00111111110010110000010100011001;
assign x[4045]= 32'b00111111110011010000010100000000;
assign x[4046]= 32'b00111111110011110000010011100111;
assign x[4047]= 32'b00111111110100010000010011001110;
assign x[4048]= 32'b00111111110100110000010010110101;
assign x[4049]= 32'b00111111110101010000010010011100;
assign x[4050]= 32'b00111111110101110000010010000011;
assign x[4051]= 32'b00111111110110000000010001101010;
assign x[4052]= 32'b00111111110110100000010001010001;
assign x[4053]= 32'b00111111110111000000010000110111;
assign x[4054]= 32'b00111111110111100000010000011110;
assign x[4055]= 32'b00111111110111110000010000000101;
assign x[4056]= 32'b00111111111000010000001111101100;
assign x[4057]= 32'b00111111111000100000001111010011;
assign x[4058]= 32'b00111111111001000000001110111010;
assign x[4059]= 32'b00111111111001010000001110100001;
assign x[4060]= 32'b00111111111001110000001110001000;
assign x[4061]= 32'b00111111111010000000001101101111;
assign x[4062]= 32'b00111111111010010000001101010110;
assign x[4063]= 32'b00111111111010110000001100111101;
assign x[4064]= 32'b00111111111011000000001100100011;
assign x[4065]= 32'b00111111111011010000001100001010;
assign x[4066]= 32'b00111111111011100000001011110001;
assign x[4067]= 32'b00111111111011110000001011011000;
assign x[4068]= 32'b00111111111100000000001010111111;
assign x[4069]= 32'b00111111111100010000001010100110;
assign x[4070]= 32'b00111111111100100000001010001101;
assign x[4071]= 32'b00111111111100110000001001110100;
assign x[4072]= 32'b00111111111101000000001001011011;
assign x[4073]= 32'b00111111111101010000001001000001;
assign x[4074]= 32'b00111111111101100000001000101000;
assign x[4075]= 32'b00111111111101110000001000001111;
assign x[4076]= 32'b00111111111110000000000111110110;
assign x[4077]= 32'b00111111111110010000000111011101;
assign x[4078]= 32'b00111111111110010000000111000100;
assign x[4079]= 32'b00111111111110100000000110101011;
assign x[4080]= 32'b00111111111110110000000110010010;
assign x[4081]= 32'b00111111111110110000000101111000;
assign x[4082]= 32'b00111111111111000000000101011111;
assign x[4083]= 32'b00111111111111000000000101000110;
assign x[4084]= 32'b00111111111111010000000100101101;
assign x[4085]= 32'b00111111111111010000000100010100;
assign x[4086]= 32'b00111111111111100000000011111011;
assign x[4087]= 32'b00111111111111100000000011100010;
assign x[4088]= 32'b00111111111111100000000011001001;
assign x[4089]= 32'b00111111111111110000000010101111;
assign x[4090]= 32'b00111111111111110000000010010110;
assign x[4091]= 32'b00111111111111110000000001111101;
assign x[4092]= 32'b00111111111111110000000001100100;
assign x[4093]= 32'b00111111111111110000000001001011;
assign x[4094]= 32'b00111111111111110000000000110010;
assign x[4095]= 32'b00111111111111110000000000011001;

    always @(posedge clk) begin
        x1_re            <=  x[address1][31:16];
        x1_im            <=  x[address1][15:0] ;
        x2_re            <=  x[address2][31:16];
        x2_im            <=  x[address2][15:0] ;
        x3_re            <=  x[address3][31:16];
        x3_im            <=  x[address3][15:0] ;
        x4_re            <=  x[address4][31:16];
        x4_im            <=  x[address4][15:0] ;
        x5_re            <=  x[address5][31:16];
        x5_im            <=  x[address5][15:0] ;
        x6_re            <=  x[address6][31:16];
        x6_im            <=  x[address6][15:0] ;
        x7_re            <=  x[address7][31:16];
        x7_im            <=  x[address7][15:0] ;
    end

endmodule
